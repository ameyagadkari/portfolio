--sync.vhd
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.game.all;

entity sync is
	port(clk_s:in std_logic;
			r_shift,l_shift,start,resetgame,pause:in std_logic;
			level_select:in std_logic_vector(2 downto 0);
			hsync,vsync:out std_logic;
			r,g,b:out std_logic_vector(3 downto 0));
end sync;

architecture sync_arch of sync is
	
	signal notstarted:std_logic:='1';--to check if game is not yet started and to display welcome message	
	signal hpos:integer range 1 to 800:=1;--pixel position including fp, bp and hsync
	signal vpos:integer range 1 to 525:=1;--pixel position including fp,bp and vsync
	signal hpos_scr:integer range 1 to 640:=1;--cursor position on screen
	signal vpos_scr:integer range 1 to 480:=1;--cursor position on screen
	signal r_bat,g_bat,b_bat,r_ball,g_ball,b_ball,r_gameover,g_gameover,b_gameover,r_lives,b_lives,g_lives,r_welmes,g_welmes,b_welmes,r_winmes,g_winmes,b_winmes,r_paused,g_paused,b_paused:std_logic_vector(3 downto 0);--rgb signals
	signal draw_bat:std_logic;	--validity signals
	signal isalive:integer:=3;--to check if lives are over
	
	signal bat_x:integer:=275; --starting x coordinate for bat
	signal bat_y:integer:=460;	--y coordinate of bat is fixed

	signal ball_x:integer:=299;--starting coordinates for ball
	signal ball_y:integer:=450;
	
	signal lives_x:integer:=550;--fixed coordinates to display lives
	signal lives_y:integer:=0;
	
	signal welmes_x:integer:=72;--fixed coordinates to display welcome message
	signal welmes_y:integer:=45;
	
	signal gameover_x:integer:=84;--fixed coordinates to display gameover
	signal gameover_y:integer:=195;
	
	signal winmes_x:integer:=90;--fixed coordinates to display winning message
	signal winmes_y:integer:=175;
	
	signal paused_x:integer:=128;--fixed coordinates to display paused message
	signal paused_y:integer:=202;
	
	signal rand_x:integer range 26 to 611:=26;--used to randomly assign x cood to bat and ball;
	signal stopball:std_logic:='0';--to stop the ball after gameover or game has been won
	
	signal l2notstarted,l3notstarted,l4notstarted,l5notstarted:std_logic:='1';--to reposition bat,ball and give initial velocity to ball at start of each level except 1st 
	signal l1complete,l2complete,l3complete,l4complete,l5complete:std_logic:='0';--to say that level is completed
	signal level_selected:std_logic:='0';--to select level at start of the game
	
	type rom_lives is array (24 downto 0)of std_logic_vector(91 downto 0);-- ROM definition of lives
	signal lives_row,lives_col: integer;--signals required by lives ROM
	signal lives_single_row: std_logic_vector(91 downto 0);
	signal lives_validity_bit: std_logic;
	
	type rom_gameover is array (89 downto 0)of std_logic_vector(471 downto 0);--ROM definition of gameover
	signal gameover_row,gameover_col: integer;--signals required by gameover ROM
	signal gameover_single_row: std_logic_vector(471 downto 0);
	signal gameover_validity_bit: std_logic;
	
	type rom_welmes is array (389 downto 0)of std_logic_vector(495 downto 0);--ROM definition of welcome message
	signal welmes_row,welmes_col: integer;--signals required by welcome ROM
	signal welmes_single_row: std_logic_vector(495 downto 0);
	signal welmes_validity_bit: std_logic;
	
	type rom_paused is array (75 downto 0)of std_logic_vector(383 downto 0);--ROM definition of pause message
	signal paused_row,paused_col: integer;--signals required by pause ROM
	signal paused_single_row: std_logic_vector(383 downto 0);
	signal paused_validity_bit: std_logic;
	
	type rom_winmes is array (129 downto 0)of std_logic_vector(459 downto 0);--ROM definition of winning message
	signal winmes_row,winmes_col: integer;--signals required by win ROM
	signal winmes_single_row: std_logic_vector(459 downto 0);
	signal winmes_validity_bit: std_logic;
	
	type rom_ball is array (12 downto 0)of std_logic_vector(12 downto 0);-- ROM definition of ball
	signal ball_row,ball_col: integer;--signals required by ball ROM
	signal ball_single_row: std_logic_vector(12 downto 0);
	signal ball_validity_bit: std_logic;
	
	signal ball_x_vel:std_logic:='1';--used to change ball movements in x and y direction after hitting a wall or brick
	signal ball_y_vel:std_logic:='0';
	signal ball_x_vel_rand:std_logic:='0';
	
	type brick_cood is array (71 downto 0) of integer;--array to store coordinates of bricks
	type brick_color is array (71 downto 0) of std_logic_vector(3 downto 0);--array to give color to each brick
	
	signal x_cood_l1:brick_cood:=--x coordinates of bricks in level1
	(20,100,180,260,340,420,500,580,
	20,100,180,260,340,420,500,580,
	20,100,180,260,340,420,500,580,
	20,100,180,260,340,420,500,580,
	20,100,180,260,340,420,500,580,
	20,100,180,260,340,420,500,580,
	20,100,180,260,340,420,500,580,
	20,100,180,260,340,420,500,580,
	20,100,180,260,340,420,500,580);
	
	signal y_cood_l1:brick_cood:=--y coordinates of bricks in level1
	(25,25,25,25,25,25,25,25,
	65,65,65,65,65,65,65,65,
	105,105,105,105,105,105,105,105,
	145,145,145,145,145,145,145,145,
	185,185,185,185,185,185,185,185,
	225,225,225,225,225,225,225,225,
	265,265,265,265,265,265,265,265,
	305,305,305,305,305,305,305,305,
	345,345,345,345,345,345,345,345);
	
	signal x_cood_l2:brick_cood:=--x coordinates of bricks in level2
	(40,80,120,160,200,240,280,
	560,520,480,440,400,360,320,
	280,240,200,160,120,80,40,
	320,360,400,440,480,520,560,others=>0);
	
	signal y_cood_l2:brick_cood:=--y coordinates of bricks in level2
	(40,60,80,100,120,140,160,
	40,60,80,100,120,140,160,
	180,200,220,240,260,280,300,
	180,200,220,240,260,280,300,others=>0);
	
	signal x_cood_l3:brick_cood:=--x coordinates of bricks in level3
	(300,260,220,180,140,100,60,20,
	340,380,420,460,500,540,580,
	300,260,220,180,140,100,60,20,
	340,380,420,460,500,540,580,
	300,260,220,180,140,100,
	340,380,420,460,500,
	300,260,220,180,140,100,
	340,380,420,460,500,
	300,260,220,180,
	340,380,420,
	300,260,220,180,
	340,380,420,
	300,260,
	340,
	300,260,
	340);
	
	signal y_cood_l3:brick_cood:=--y coordinates of bricks in level3
	(25,45,65,85,105,125,145,165,
	45,65,85,105,125,145,165,
	325,305,285,265,245,225,205,185,
	305,285,265,245,225,205,185,
	65,85,105,125,145,165,
	85,105,125,145,165,
	285,265,245,225,205,185,
	265,245,225,205,185,
	105,125,145,165,
	125,145,165,
	245,225,205,185,
	225,205,185,
	145,165,
	165,
	205,185,
	185);
	
	signal x_cood_l4:brick_cood:=--x coordinates of bricks in level4
	(40,80,120,160,200,240,280,
	560,520,480,440,400,360,320,
	280,240,200,160,120,80,40,
	320,360,400,440,480,520,560,
	40,40,40,40,40,40,40,40,40,
	560,560,560,560,560,560,560,560,560,
	100,150,200,250,300,350,400,450,500,
	100,150,200,250,300,350,400,450,500,others=>0);
	
	signal y_cood_l4:brick_cood:=--y coordinates of bricks in level4
	(40,60,80,100,120,140,160,
	40,60,80,100,120,140,160,
	180,200,220,240,260,280,300,
	180,200,220,240,260,280,300,
	70,95,120,145,170,195,220,245,270,
	70,95,120,145,170,195,220,245,270,
	40,40,40,40,40,40,40,40,40,
	300,300,300,300,300,300,300,300,300,others=>0);
	
	signal x_cood_l5:brick_cood:=--x coordinates of bricks in level5
	(20,60,100,140,180,220,260,
	340,380,420,460,500,540,580,
	140,140,140,140,140,140,140,140,140,140,140,
	460,460,460,460,460,460,460,460,460,460,460,others=>0);
	
	signal y_cood_l5:brick_cood:=--y coordinates of bricks in level5
	(85,65,45,25,45,65,85,
	85,65,45,25,45,65,85,
	65,90,115,140,165,190,215,240,265,290,315,
	65,90,115,140,165,190,215,240,265,290,315,others=>0);
	
	
	signal is_destroyed_l1,coll_x_l1,coll_y_l1,draw_l1:std_logic_vector(71 downto 0):=x"000000000000000000";--for level 1
	signal is_destroyed_l2,coll_x_l2,coll_y_l2,draw_l2:std_logic_vector(71 downto 44):=x"0000000";--for level 2
	signal is_destroyed_l3,coll_x_l3,coll_y_l3,draw_l3:std_logic_vector(71 downto 0):=x"000000000000000000";--for level 3
	signal is_destroyed_l4,coll_x_l4,coll_y_l4,draw_l4:std_logic_vector(71 downto 8):=x"0000000000000000";--for level 4
	signal is_destroyed_l5,coll_x_l5,coll_y_l5,draw_l5:std_logic_vector(71 downto 36):=x"000000000";--for level 5
	
	signal r_brick,g_brick,b_brick:brick_color;--rgb for bricks

	constant lives0_rom: rom_lives:= --lives 0 image
	(
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"000780f0038747c020f3ffe",
x"0018c318038cc9e07073078",
x"0018c318038c40e07072078",
x"0038e71c000e00707872078",
x"0038e71c000f0070b870078",
x"0038e71c0007cff0b870078",
x"0038e71c0003cc711c70078",
x"0038e71c0388cc611c70078",
x"0038e71c038cc6e31e70078",
x"0038e71c038b8387bf70078",
x"0038e71c000000000000078",
x"0018c318000000000060078",
x"0018c318000000000070078",
x"000780f00000000000601fe",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000"
);

	constant lives1_rom: rom_lives:= --lives 1 image
	(
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"001fc0f0038747c020f3ffe",
x"00070318038cc9e07073078",
x"00070318038c40e07072078",
x"0007071c000e00707872078",
x"0007071c000f0070b870078",
x"0007071c0007cff0b870078",
x"0007071c0003cc711c70078",
x"0007071c0388cc611c70078",
x"0007071c038cc6e31e70078",
x"0007071c038b8387bf70078",
x"0007071c000000000000078",
x"0007c318000000000060078",
x"00078318000000000070078",
x"000600f00000000000601fe",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000"
);

	constant lives2_rom: rom_lives:= --lives 2 image
	(
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"001fe0f0038747c020f3ffe",
x"001fc318038cc9e07073078",
x"003fc318038c40e07072078",
x"0020871c000e00707872078",
x"0001071c000f0070b870078",
x"0002071c0007cff0b870078",
x"0006071c0003cc711c70078",
x"000c071c0388cc611c70078",
x"001c071c038cc6e31e70078",
x"001c071c038b8387bf70078",
x"001c071c000000000000078",
x"001e2318000000000060078",
x"000fc318000000000070078",
x"000780f00000000000601fe",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000"
);

	constant lives3_rom: rom_lives := --lives 3 image
	(
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"0007e0f0038747c020f3ffe",
x"0008f318038cc9e07073078",
x"00186318038c40e07072078",
x"0038071c000e00707872078",
x"0038071c000f0070b870078",
x"003c071c0007cff0b870078",
x"003e071c0003cc711c70078",
x"001f871c0388cc611c70078",
x"0006071c038cc6e31e70078",
x"001c071c038b8387bf70078",
x"001c071c000000000000078",
x"001e2318000000000060078",
x"001fc318000000000070078",
x"000f80f00000000000601fe",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000",
x"00000000000000000000000"
);


	constant winmes_rom: rom_winmes:= --winning image
(
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000780000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000fc0000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000000000000000000000013c0000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000000000000000000000013c0000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000002380000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000006000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000",
x"008003fcffefff83fe00ff800fff83fe0001fff81fff07fcfffffc00fff80007e00f000001fc004000f81fff1ffe0007cc1f303e001ff003ffe",
x"00c000f03f83fc007807fff003fc007800003f8007f800f0fffff0001fe0001e781f800007ff00e003fe07fc07f0000e3c38f0ff800fc0007f8",
x"00e000603f81fc00301f81f801fc003000003f8003f80060f80fe0000fc0003c3c27c0001fff00e0063f03fc03f0001c1c70718fc007c0003f0",
x"00f000601f80fc00203f007e00fc002000001f8001f80040e007e0000fc0007c3c07c0003c3f01f0001f81fc03f0003c0cf03007e007c0003f0",
x"00f800601f80fe00603f003f00fe006000001f8001fc00c0c007e0000fc0007c3e07c000381f01f0080f80fe03f0003e04f81203e007c0003f0",
x"00f800601f80fe00403f003f80fe004000001f8001fc0080c007e0000fc0007c3e07c000780701f8000f807f03f0003f00fc0003e007c0003f0",
x"00fc00601f807e00c03f001f807e00c000001f8000fc01818007e0000fc000fc3f07c000700003f8000fc07f83f0003fc0ff0003f007c0003f0",
x"00fe00601f807fffc03f001fc07fffc000001f8000ffff818007e0000fc000f83f07c000f80002fc0007c03f83f0001fe07f8001f007c0003f0",
x"00ff00601f803fff803f000fc03fff8000001f80007fff010007e0000fc000f83f07c000f80006fc0007c01fc3f0001ff07fc001f007c0003f0",
x"00ff80601f803f81807f800fc03f818000001f80007f03000007e0000fc000f83f07c000f800047c0fffc00fe3f0000ff83fe3fff007c0003f0",
x"00ffc0601f801f8101ffe00fc01f810000003f80003f02000007e0000fc000f83f07c000fc00047e0f07c007f3f00003f80fe3c1f007c0003f0",
x"00dfc0601f801f830000000fe01f830000003fc0003f06000007e003ffc0007c3e07c000ff00083e0f078007fff00001fc07f3c1e00fc00fff0",
x"00dfe0601f801fc20000000fe01fc20000006fc0003f84000007e01fffc0007c3e07c0007fc0083f0f078003fff000107c41f3c1e30fc07fff0",
x"00cff0601f800fc60000000fc00fc60000004fe0001f8c000007e03f8fc0007c3c07c0003ff0181f070f0001fff000183860e1c3c78fc0fe3f0",
x"00c7f8601f800fe60000000fc00fe6000000c7e0001fcc000007e07e0fc0003c3c07c0001fc0181f878f0000f3f0001c3870e1e3c7d7c1f83f0",
x"00c3fc601f8007ec0000000fc007ec00000187f0000fd8000007e07e0fc0001e787ff8000f00381fc39e0000e3f0001e3078c0e787e7c1f83f0",
x"00c1fe601f8007fc0000001fc007fc00000183f0000ff8000007e0fc0fc00007e07fe0001e007e3fe0f8000183f00013e04f803e03c7f3f03f0",
x"00c0fe601f8003f80020001f8003f800000301f80007f0000007e0fc0fc000000007c0003e0000000000000303f0000000000000000003f03f0",
x"00c0ff601f8003f80030001f8003f800000201fc0007f0000007e0fc0fc00000000780003e0000000000000603f0000000000000000003f03f0",
x"00c07fe01f8003f00030003f0003f000000600fc0007e0000007e0fc0fc00000000700003e0000000000001c03f0000000000000000003f03f0",
x"00c03fe01f8001f00038003e0001f000000c00fe0003e0000007e0fe0fc00000000600007e0200000000003803f0000000000000000003f83f0",
x"00c01fe01f8001f0003e007c0001f000000c007e0003e0000007e07e0fc00000000600003f0600000000006003f0000000000000000001f83f0",
x"00c00fe03f8000e0003f81f80000e000001c007f0001c0000007e03f8fc00000000400003ffc0000000001e003f0000000000000000000fe3f0",
x"01e00ff83f8000e00033ffe00000e000003c007f8001c000000ff01fffe00000000000001ff80000000003e007f00000000000000000007fff8",
x"07f807feffe0004000207f8000004000007f01ffe0008000007ffc07fff800000000000007e0000000000ff81ffe0000000000000000001fffe",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"001fffff7ffe0c0ff7ffc1ff007fc000001f01ff7fc3c00008003fc007fc00001000c000001f0001001e0f0fffbffe003f9f800fc001fff8000",
x"003ffff80ff00c03c1fe003c03fff800007fc07c3f07e0000c000f001fff00003800c000007fc003807f7f83fc07f8000fffc03cf0003f80000",
x"003e03f807e00e0180fe00180fc0fc0000c7e07c1f09f0000e0006007e0fc0003801c00000c7e003801f9f81f803f0000fe7c07878003f80000",
x"003801f807e01e01807e00101f803f000003f07c1f01f0000f000600fc07e0003801e0000003f007c01f0f81f803f0000fc3e0f878001f80000",
x"003001f807e01f01807f00301f801f800101f07c1f01f0000f800601f803f0007c03e0000101f007c01f0f81f803f0000f83e0f87c001f80000",
x"002001f807e03f01807f00201f801fc00001f07c1f01f0000f800603f001f8007c03f0000001f007c01f0f81f803f0000f83e0f87c001f80000",
x"002041f807e03f81803f00601f800fc00001f87c1f01f0000fc00603f001f800fc03f0000001f80fe01f0f01f803f0000f83e1f87e001f80000",
x"002041f807e07f81803fffe01f800fe00000f87c1f01f0000fe00607e001fc00fe07f0000000f80be01f1c01f803f0000f83e1f07e001f80000",
x"000041f807e07fc1801fffc01f8007e00000f87c1f01f0000ff00607e000fc00fe07f8000000f813f01f3801f803f0000f83e1f07e001f80000",
x"000041f807e05fc1801fc0c03fc007e001fff87c1f01f0000ff80607e000fc01ff0df80001fff813f01fe001f803f0000f83e1f07e001f80000",
x"000061f807e0cfe1800fc080fff007e001e0f87c1f01f0000ffc060fe000fc01bf0dfc0001e0f831f81f0f01f803f0000f83e1f07e003f80000",
x"000071f807e08fe1800fc180000007f001e0f07c1f01f0000dfc060fe000fe013f08fc0001e0f021f81f0f81f803f0000f83e0f87c003fc0000",
x"00007ff807e187e1800fe100000007f001e0f07c1f01f0000dfe060fe000fe031f98fc0001e0f060f81f0f81fffff0000f83e0f87c006fc0000",
x"00007ff807e107f18007e300000007e000e1e07c3f01f0000cff060fe000fe021f907e0000e1e040fc1f0f81fffff0000f83e0f878004fe0000",
x"000071f807e303f18007f300000007e000f1e07e7f01f0000c7f860fe000fc061fb07e0000f1e0c07c1f0701f803f0000f83e0787800c7e0000",
x"000061f807e303f98003f600000007e00073c03fdf1ffe000c3fc607e000fc060ff07f000073c0c0fe0f8e01f803f0000fc3e03cf00187f0000",
x"000041f807e603f98003fe0000000fe0001f001f1f1ff8000c1fe607e000fc040fe03f00001f01f1ff03f801f803f0000fe3f80fc00183f0000",
x"001041f807e601fd8001fc0010000fc0000000001f01f0000c0fe607e001fc0c0fe03f000000000000000001f803f00000000000000301f8000",
x"001841f807e401fd8001fc0018000fc0000000001f01e0000c0ff603f001f80c07e01f800000000000000001f803f00000000000000201fc000",
x"001841f807ec00ff8001f80018001f80000000001f01c0000c07fe03f001f80807e01f800000000000000001f803f00000000000000600fc000",
x"001801f807fc00ff8000f8001c001f00000000001f0180000c03fe01f803f01803f01fc00000000000000001f803f00000000000000c00fe000",
x"001c01f807f8007f8000f8001f003e00000000001f0180000c01fe00f807e01003f00fc00000000000000001f803f00000000000000c007e000",
x"001f01f807f8007f800070001fc0fc00000000001f0100000c00fe007e0fc03003f80fe00000000000000001f803f00000000000001c007f000",
x"001ffff80ff0007f8000700019fff000000000001f0000001e00ff803fff003803fc0fe00000000000000003fc07f80000000000003c007f800",
x"001fffff7ff0003ff0002000103fc000000000001fc000007f807fe007fc00fe0fff3ff8000000000000000fffbffe0000000000007f01ffe00",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000003f0403ffe07ffc1ffff07ffc00ff80008003fc007fc0000ff00000000000000000000000000000000",
x"0000000000000000000000000000000000ffc4007f001fe003c7f80ff007fff000c000f001fff0003ffe0000000000000000000000000000000",
x"0000000000000000000000000000000001e0fc007f000fe00183f807e01f81f800e0006007e0fc00f03f8000000000000000000000000000000",
x"0000000000000000000000000000000003c03c003f0007e00101fc07e03f007e00f000600fc07e01c00fc000000000000000000000000000000",
x"0000000000000000000000000000000007801c003f0007f00300fe07e03f003f00f800601f803f030007e000000000000000000000000000000",
x"0000000000000000000000000000000007800c003f0007f002007e07e03f003f80f800603f001f820007f000000000000000000000000000000",
x"00000000000000000000000000000000078004003f0003f006007f07e03f001f80fc00603f001f800003f000000000000000000000000000000",
x"0000000000000000000000000000000007c004003f0003fffe003f87e03f001fc0fe00607e001fc00003f800000000000000000000000000000",
x"0000000000000000000000000000000007e004003f0001fffc001fc7e03f000fc0ff00607e000fc00003f800000000000000000000000000000",
x"0000000000000000000000000000000007f800003f0001fc0c001fc7e07f800fc0ff80607e000fc00001f800000000000000000000000000000",
x"0000000000000000000000000000000007fe00003f0000fc08000fe7e1ffe00fc0ffc060fe000fc00001f800000000000000000000000000000",
x"0000000000000000000000000000000003ff80003f0000fc180007ffe000000fe0dfc060fe000fe00001fc00000000000000000000000000000",
x"0000000000000000000000000000000001ffe0003f0000fe10001fffe000000fe0dfe060fe000fe00001fc00000000000000000000000000000",
x"0000000000000000000000000000000000fff0003f00007e30007f07e000000fc0cff060fe000fe00001f800000000000000000000000000000",
x"00000000000000000000000000000000003ff8003f00007f30007e07e000000fc0c7f860fe000fc00001f800000000000000000000000000000",
x"00000000000000000000000000000000000ff8003f00003f6000fc07e000000fc0c3fc607e000fc00001f800000000000000000000000000000",
x"000000000000000000000000000000000001fc003f00003fe000fc07e000001fc0c1fe607e000fc00003f800000000000000000000000000000",
x"000000000000000000000000000000000200fc003f00001fc001f807e020001f80c0fe607e001fc20003f000000000000000000000000000000",
x"0000000000000000000000000000000002007c403f01001fc001fc07e030001f80c0ff603f001f820003f000000000000000000000000000000",
x"0000000000000000000000000000000003003c403f01001f8000fc07e030003f00c07fe03f001f830007e000000000000000000000000000000",
x"0000000000000000000000000000000003003c603f03000f8000fc07e038003e00c03fe01f803f03000fc000000000000000000000000000000",
x"0000000000000000000000000000000003c038703f07000f8000fe07e03e007c00c01fe00f807e03c01f8000000000000000000000000000000",
x"0000000000000000000000000000000003e0f0783f0f000700007f07e03f81f800c00fe007e0fc03f07f0000000000000000000000000000000",
x"00000000000000000000000000000000027fe07fffff000700003ffff033ffe001e00ff803fff0023ffc0000000000000000000000000000000",
x"00000000000000000000000000000000021f807fffff0002000007fffc207f8007f807fe007fc0020ff00000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"

);
	constant gameover_rom: rom_gameover:= --gameover image
(
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000000000000000000000000f0000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000000000000000000000001f8000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000278000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000278000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000470000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000400000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000c00000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000800000000000000000000000000000000000000",
x"0010007f9ffdfff07fc01ff001fff07fc0003fff03ffe0ff9fffff801fff0000fc01e000003f8008001f03ffe3ffc000f983e607c003fe007ffc00",
x"0018001e07f07f800f00fffe007f800f000007f000ff001e1ffffe0003fc0003cf03f00000ffe01c007fc0ff80fe0001c7871e1ff001f8000ff000",
x"001c000c07f03f800603f03f003f8006000007f0007f000c1f01fc0001f800078784f80003ffe01c00c7e07f807e0003838e0e31f800f80007e000",
x"001e000c03f01f800407e00fc01f8004000003f0003f00081c00fc0001f8000f8780f8000787e03e0003f03f807e0007819e0600fc00f80007e000",
x"001f000c03f01fc00c07e007e01fc00c000003f0003f80181800fc0001f8000f87c0f8000703e03e0101f01fc07e0007c09f02407c00f80007e000",
x"001f000c03f01fc00807e007f01fc008000003f0003f80101800fc0001f8000f87c0f8000f00e03f0001f00fe07e0007e01f80007c00f80007e000",
x"001f800c03f00fc01807e003f00fc018000003f0001f80303000fc0001f8001f87e0f8000e00007f0001f80ff07e0007f81fe0007e00f80007e000",
x"001fc00c03f00ffff807e003f80ffff8000003f0001ffff03000fc0001f8001f07e0f8001f00005f8000f807f07e0003fc0ff0003e00f80007e000",
x"001fe00c03f007fff007e001f807fff0000003f0000fffe02000fc0001f8001f07e0f8001f0000df8000f803f87e0003fe0ff8003e00f80007e000",
x"001ff00c03f007f0300ff001f807f030000003f0000fe0600000fc0001f8001f07e0f8001f00008f81fff801fc7e0001ff07fc7ffe00f80007e000",
x"001ff80c03f003f0203ffc01f803f020000007f00007e0400000fc0001f8001f07e0f8001f80008fc1e0f800fe7e00007f01fc783e00f80007e000",
x"001bf80c03f003f060000001fc03f060000007f80007e0c00000fc007ff8000f87c0f8001fe00107c1e0f000fffe00003f80fe783c01f801ffe000",
x"001bfc0c03f003f840000001fc03f84000000df80007f0800000fc03fff8000f87c0f8000ff80107e1e0f0007ffe00020f883e783c61f80fffe000",
x"0019fe0c03f001f8c0000001f801f8c0000009fc0003f1800000fc07f1f8000f8780f80007fe0303e0e1e0003ffe0003070c1c3878f1f81fc7e000",
x"0018ff0c03f001fcc0000001f801fcc0000018fc0003f9800000fc0fc1f800078780f80003f80303f0f1e0001e7e0003870e1c3c78faf83f07e000",
x"00187f8c03f000fd80000001f800fd80000030fe0001fb000000fc0fc1f80003cf0fff0001e00703f873c0001c7e0003c60f181cf0fcf83f07e000",
x"00183fcc03f000ff80000003f800ff800000307e0001ff000000fc1f81f80000fc0ffc0003c00fc7fc1f0000307e00027c09f007c078fe7e07e000",
x"00181fcc03f0007f00040003f0007f000000603f0000fe000000fc1f81f800000000f80007c0000000000000607e0000000000000000007e07e000",
x"00181fec03f0007f00060003f0007f000000403f8000fe000000fc1f81f800000000f00007c0000000000000c07e0000000000000000007e07e000",
x"00180ffc03f0007e00060007e0007e000000c01f8000fc000000fc1f81f800000000e00007c0000000000003807e0000000000000000007e07e000",
x"001807fc03f0003e00070007c0003e000001801fc0007c000000fc1fc1f800000000c0000fc0400000000007007e0000000000000000007f07e000",
x"001803fc03f0003e0007c00f80003e000001800fc0007c000000fc0fc1f800000000c00007e0c0000000000c007e0000000000000000003f07e000",
x"001801fc07f0001c0007f03f00001c000003800fe00038000000fc07f1f800000000800007ff80000000003c007e0000000000000000001fc7e000",
x"003c01ff07f0001c00067ffc00001c000007800ff00038000001fe03fffc00000000000003ff00000000007c00fe0000000000000000000ffff000",
x"00ff00ffdffc000800040ff000000800000fe03ffc001000000fff80ffff00000000000000fc0000000001ff03ffc0000000000000000003fffc00",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000380700e1fe0fff87ffffc000c00000ff8003ffffefffc181fefff83fe00ff8000e01c0380000000000000000000000000",
x"0000000000000000000007c0f81f0ff01fe0ffffe0000c00003ffe007ffff01fe0180783fc007807fff001f03e07c0000000000000000000000000",
x"000000000000000000000fe1fc3f87f00fc0f80fe0001e0000fc1f807c07f00fc01c0301fc00301f81f803f87f0fe0000000000000000000000000",
x"0000000000000000000007c0f81f03f80fc0e007e0001e0001f80fc07003f00fc03c0300fc00203f007e01f03e07c0000000000000000000000000",
x"000000000000000000000380700e01fc0fc0c007e0003e0003f007e06003f00fc03e0300fe00603f003f00e01c0380000000000000000000000000",
x"000000000000000000000000000000fc0fc08007e0003f0007e003f04003f00fc07e0300fe00403f003f8000000000000000000000000000000000",
x"000000000000000000000000000000fe0fc08107e0007f0007e003f04083f00fc07f03007e00c03f001f8000000000000000000000000000000000",
x"0000000000000000000000000000007f0fc08107e0007f800fc003f84083f00fc0ff03007fffc03f001fc000000000000000000000000000000000",
x"0000000000000000000001002004003f8fc00107e0005f800fc001f80083f00fc0ff83003fff803f000fc040080100000000000000000000000000",
x"0000000000000000000001002004003f8fc00107e000df800fc001f80083f00fc0bf83003f81807f800fc040080100000000000000000000000000",
x"0000000000000000000001002004001fcfc00187e0008fc01fc001f800c3f00fc19fc3001f8101ffe00fc040080100000000000000000000000000",
x"0000000000000000000001002004000fffc001c7e0018fc01fc001fc00e3f00fc11fc3001f830000000fe040080100000000000000000000000000",
x"000000000000000000000380700e003fffc001ffe00107e01fc001fc00fff00fc30fc3001fc20000000fe0e01c0380000000000000000000000000",
x"000000000000000000000380700e00fe0fc001ffe00307e01fc001fc00fff00fc20fe3000fc60000000fc0e01c0380000000000000000000000000",
x"000000000000000000000380700e00fc0fc001c7e00307f01fc001f800e3f00fc607e3000fe60000000fc0e01c0380000000000000000000000000",
x"000000000000000000000380700e01f80fc00187e00603f00fc001f800c3f00fc607f30007ec0000000fc0e01c0380000000000000000000000000",
x"0000000000000000000007c0f81f01f80fc00107e00603f00fc001f80083f00fcc07f30007fc0000001fc1f03e07c0000000000000000000000000",
x"0000000000000000000007c0f81f03f00fc04107e00401f80fc003f82083f00fcc03fb0003f80020001f81f03e07c0000000000000000000000000",
x"0000000000000000000007c0f81f03f80fc06107e00c01f807e003f03083f00fc803fb0003f80030001f81f03e07c0000000000000000000000000",
x"0000000000000000000007c0f81f01f80fc06107e00801fc07e003f03083f00fd801ff0003f00030003f01f03e07c0000000000000000000000000",
x"0000000000000000000007c0f81f01f80fc06007e01800fc03f007e03003f00ff801ff0001f00038003e01f03e07c0000000000000000000000000",
x"000000000000000000000fe1fc3f81fc0fc07007e01800fe01f00fc03803f00ff000ff0001f0003e007c03f87f0fe0000000000000000000000000",
x"000000000000000000000fe1fc3f80fe0fc07c07e030007e00fc1f803e03f00ff000ff0000e0003f81f803f87f0fe0000000000000000000000000",
x"0000000000000000000007c0f81f007fffe07fffe078007f007ffe003ffff01fe000ff0000e00033ffe001f03e07c0000000000000000000000000",
x"000000000000000000000380700e000ffff87ffffdff03ffc00ff8003ffffeffe0007fe0004000207f8000e01c0380000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
);

	constant welmes_rom: rom_welmes:= --welcome message image
(
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000078000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000fc000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000013c000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000013c000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000238000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000600000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000400000000000000000000000000000000000000000",
x"000000000000000000000000000000000001e001000c0000fc103c01f003e67f3f00f078007ffc01804003c1e3fe007ffc00000000000000000000000000",
x"00000000000000000000000000000000001f8003800c0003ff107e07fc071e1fff83fbfc000ff00380e00feff0fc000ff000000000000000000000000000",
x"00000000000000000000000000000000007c0003801c000783f07e0c7e0e0e1fcf80fcfc0007e00300e003f3f0f80007e000000000000000000000000000",
x"0000000000000000000000000000000000f80003801e000f00f07e003f1e061f87c0f87c0007e00301f003e1f0f80007e000000000000000000000000000",
x"0000000000000000000000000000000001f00007c03e001e00703c101f1f021f07c0f87c0007e00701f003e1f0f80007e000000000000000000000000000",
x"0000000000000000000000000000000003e00007c03f001e003000001f1f801f07c0f87c0007e00601f803e1f0f80007e000000000000000000000000000",
x"0000000000000000000000000000000007c0000fc03f001e001000001f9fe01f07c0f8780007e00603f803e1e0f80007e000000000000000000000000000",
x"000000000000000000000000000000000f80000fe07f001f001000000f8ff01f07c0f8e00007e00e02fc03e380f80007e000000000000000000000000000",
x"000000000000000000000000000000000f80000fe07f801f801000000f8ff81f07c0f9c00007e00c06fc03e700f80007e000000000000000000000000000",
x"000000000000000000000000000000001f80001ff0df801fe000001fff87fc1f07c0ff000007e00c047c03fc00f80007e000000000000000000000000000",
x"000000000000000000000000000000001ffe001bf0dfc01ff800001e0f81fc1f07c0f8780007e00c047e03e1e0f80007e000000000000000000000000000",
x"000000000000000000000000000000001f1f0013f08fc00ffe00001e0f00fe1f07c0f87c01ffe01c083e03e1f0f801ffe000000000000000000000000000",
x"000000000000000000000000000000001f0f8031f98fc007ff803c1e0f083e1f07c0f87c0fffe018083f03e1f0f80fffe000000000000000000000000000",
x"000000000000000000000000000000003f07c021f907e003ffc07e0e1e0c1c1f07c0f87c1fc7e018181f03e1f0f81fc7e000000000000000000000000000",
x"000000000000000000000000000000003f07c061fb07e000ffe07e0f1e0e1c1f07c0f8383f07e038181f83e0e0f83f07e000000000000000000000000000",
x"000000000000000000000000000000003f07c060ff07f0003fe07e073c0f181f87c07c703f07e030381fc1f1c0f83f07e000000000000000000000000000",
x"000000000000000000000000000000003f07e040fe03f00007f03c01f009f01fc7f01fc07e07e0307e3fe07f00f87e07e000000000000000000000000000",
x"000000000000000000000000000000001f07e0c0fe03f00803f0000000000000000000007e07e0700000000000f87e07e000000000000000000000000000",
x"000000000000000000000000000000001f07c0c07e01f80801f0000000000000000000007e07e0600000000000f87e07e000000000000000000000000000",
x"000000000000000000000000000000001f07c0807e01f80c00f0000000000000000000007e07e0600000000000f87e07e000000000000000000000000000",
x"000000000000000000000000000000000f87c1803f01fc0c00f0000000000000000000007f07e0e00000000000f87f07e000000000000000000000000000",
x"000000000000000000000000000000000f8781003f00fc0f00e0000000000000000000003f07e0c00000000000f83f07e000000000000000000000000000",
x"00000000000000000000000000000000078783003f80fe0f83c0000000000000000000001fc7e0c00000000000f81fc7e000000000000000000000000000",
x"0000000000000000000000000000000003ce03803fc0fe09ff80000000000000000000000ffff0c00000000000fc0ffff000000000000000000000000000",
x"0000000000000000000000000000000000fc0fe0fff3ff887e000000000000000000000003fffd800000000000fe03fffc00000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000060000000000000000000018000000000000000000000000000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000c0000000000000000000030000000000000000000000000000000000000000000000000000000000000000000000000000",
x"00000000000000000000000003800000000000000000000e0000000000000000000000000000000000000000000000000000000000000000000000000000",
x"00000000000000000000000003000000000000000000000c0000000000000000000000000000000000000000000000000000000000000000000000000000",
x"00000000000000000000000007000000000000000000001c0000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000600000000000000000000180000000000000000000000000000000000000000000000000000000000000000000000000000",
x"00000003e0000400300003f047e0fff8001000c0000fc11f83fff800400300003f040f01e007c007c0ff81f0007e0800ff81f00010007c03fffff0000000",
x"0000000e38000e0030000ffc47e01fc0003800c0003ff11f83fff000e0030000ffc41f83f01ff01ff03f07fc01ff88003f07fc003801ff03ffffc0000000",
x"0000001e3c000e0070001e0fc7f00f80003801c000783f1fc3ffe000e0070001e0fc1f84f821f831f83e0c7e03c1f8003e0c7e0038031f83e03f80000000",
x"0000001c1e000e0078003c03c7e00f80003801e000f00f1f83ffe000e0078003c03c1f80f840fc00fc3e003f078078003e003f007c000fc3801f80000000",
x"0000003c1e001f00f8007801c1c00f80007c03e001e0070707ffc001f00f8007801c0f00f800fc407c3e101f0f0038003e101f007c0407c3001f80000000",
x"0000003c1f001f00fc007800c0000f80007c03f001e0030006018001f00fc007800c0000f8007c007c3e001f0f0018003e001f007c0007c3001f80000000",
x"0000007c1f003f00fc00780040000f8000fc03f001e0010004030003f00fc00780040000f8007e007e3e001f8f0008003e001f80fe0007e6001f80000000",
x"0000007c1f003f81fc007c0040000f8000fe07f001f0010000060003f81fc007c0040000f8007e003e3e000f8f8008003e000f80be0003e6001f80000000",
x"0000007c1f003f81fe007e0040000f8000fe07f801f80100000e0003f81fe007e0040000f8003e003e3e000f8fc008003e000f813f0003e4001f80000000",
x"0000007c1f807fc37e007f8000000f8001ff0df801fe0000001c0007fc37e007f8000000f8003e7ffe3e1fff8ff000003e1fff813f07ffe0001f80000000",
x"000000fc1f806fc37f007fe000000f8001bf0dfc01ff800000380006fc37f007fe000000f8003e783e3e1e0f8ffc00003e1e0f831f8783e0001f80000000",
x"000000fc1f804fc23f003ff800000f80013f08fc00ffe00000780004fc23f003ff800000f8003c783c3e1e0f07ff00003e1e0f021f8783c0001f80000000",
x"000000fc1f80c7e63f001ffe00000f80031f98fc007ff8000070000c7e63f001ffe00f00f8383c783c3e1e0f03ffc0003e1e0f060f8783c0001f80000000",
x"000000fc1f8087e41f800fff00000f80021f907e003ffc0000f000087e41f800fff01f80f87c7838783e0e1e01ffe0003e0e1e040fc38780001f80000000",
x"000000fc1f8187ec1f8003ff80000f80061fb07e000ffe0001f000187ec1f8003ff81f80f87c783c783e0f1e007ff0003e0f1e0c07c3c780001f80000000",
x"0000007c1f8183fc1fc000ff80000f80060ff07f0003fe0001f000183fc1fc000ff81f8fff3cf01cf03e073c001ff0003e073c0c0fe1cf00001f80000000",
x"0000007c1f0103f80fc0001fc0000f80040fe03f00007f0001e000103f80fc0001fc0f0ffc0fc007c03e01f00003f8003e01f01f1ff07c00001f80000000",
x"0000007c1f0303f80fc0200fc0000f800c0fe03f00803f0003f000303f80fc0200fc0000f8000000003e00000401f8003e00000000000000001f80000000",
x"0000007c1f0301f807e02007c0000f800c07e01f80801f0003f008301f807e02007c0000f0000000003e00000400f8003e00000000000000001f80000000",
x"0000003c1f0201f807e03003c0000f800807e01f80c00f0003f010201f807e03003c0000e0000000003e0000060078003e00000000000000001f80000000",
x"0000003c1e0600fc07f03003c0000fc81803f01fc0c00f0003fc30600fc07f03003c0000c0000000003e0000060078003e00000000000000001f80000000",
x"0000001c1e0400fc03f03c0380000ff01003f00fc0f00e0001ffe0400fc03f03c0380000c0000000003e0000078070003e00000000000000001f80000000",
x"0000001e1c0c00fe03f83e0f00000fc03003f80fe0f83c0001ffe0c00fe03f83e0f0000080000000003e000007c1e0003e00000000000000001f80000000",
x"0000000e380e00ff03f827fe00000f003803fc0fe09ff80000ffc0e00ff03f827fe0000000000000003f000004ffc0003f00000000000000003fc0000000",
x"00000003e03f83ffcffe21f800000c00fe0fff3ff887e000003f03f83ffcffe21f80000000000000003f8000043f00003f8000000000000001fff0000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007800000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fc00000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013c00000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013c00000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000023800000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040000000000000000000000000",
x"0000000000000000001fff01fff7ffc00ff8007ffff83ffe000f00f07801ffff0001f00010003f03fff0607f83c007c0004000f81fff1ffe000000000000",
x"00000000000000000003f8007f80ff007fff001fc3fc07f8001f83fbfc07fff80007fc003800f3c07f80601e07e01c7000e003fe07fc07f0000000000000",
x"00000000000000000003f8003f007e01f81f801fc1fc03f00027c0fcfc1fe1f8000c7e003801e1e03f00700c07e03c7800e0063f03fc03f0000000000000",
x"00000000000000000001f8003f007e03f007e00fc0fe03f00007c0f87c3f81f800003f007c03e1e03f00f00c07e0383c01f0001f81fc03f0000000000000",
x"00000000000000000001f8003f007e03f003f00fc07f03f00007c0f87c3f01f800101f007c03e1f03f00f80c03c0783c01f0080f80fe03f0000000000000",
x"00000000000000000001f8003f007e03f003f80fc03f03f00007c0f87c7f01f800001f007c03e1f03f01f80c0000783e01f8000f807f03f0000000000000",
x"00000000000000000001f8003f007e03f001f80fc03f83f00007c0f8787f01f800001f80fe07e1f83f01fc0c0000f83e03f8000fc07f83f0000000000000",
x"00000000000000000001f8003f007e03f001fc0fc01fc3f00007c0f8e07f01f800000f80be07c1f83f03fc0c0000f83e02fc0007c03f83f0000000000000",
x"00000000000000000001f8003f007e03f000fc0fc00fe3f00007c0f9c07f01f800000f813f07c1f83f03fe0c0000f83e06fc0007c01fc3f0000000000000",
x"00000000000000000001f8003f007e07f800fc0fc00fe3f00007c0ff003f01f8001fff813f07c1f83f02fe0c0000f83f047c0fffc00fe3f0000000000000",
x"00000000000000000001f8003f007e1ffe00fc0fc007f3f00007c0f8781f81f8001e0f831f87c1f83f067f0c0001f83f047e0f07c007f3f0000000000000",
x"00000000000000000001f8003f007e000000fe0fc003fff00007c0f87c0fe1f8001e0f021f83e1f03f047f0c0001f83f083e0f078007fff0000000000000",
x"00000000000000000001f8003ffffe000000fe0fc00ffff00007c0f87c07fff8001e0f060f83e1f03f0c3f0c03c1f83f083f0f078003fff0000000000000",
x"00000000000000000001f8003ffffe000000fc0fc03f83f00007c0f87c01fff8000e1e040fc3e1e03f083f8c07e1f83f181f070f0001fff0000000000000",
x"00000000000000000001f8003f007e000000fc0fc03f03f00007c0f83807e1f8000f1e0c07c1e1e03f181f8c07e1f83f181f878f0000f3f0000000000000",
x"00000000000000000001f8003f007e000000fc0fc07e03f0007ff87c700fc1f800073c0c0fe0f3c03f181fcc07e0f83f381fc39e0000e3f0000000000000",
x"00000000000000000001f8003f007e000001fc0fc07e03f0007fe01fc01f81f80001f01f1ff03f003f301fcc03c0f83e7e3fe0f8000183f0000000000000",
x"00000000000000000001f8003f007e020001f80fc0fc03f00007c000003f81f800000000000000003f300fec0000f83e00000000000303f0000000000000",
x"00000000000000000201f8083f007e030001f80fc0fe03f000078000003f81f800000000000000003f200fec0000f83e00000000000603f0000000000000",
x"00000000000000000201f8083f007e030003f00fc07e03f000070000003f81f800000000000000003f6007fc0000783e00000000001c03f0000000000000",
x"00000000000000000301f8183f007e038003e00fc07e03f000060000001f81f800000000000000003fe007fc0000783c00000000003803f0000000000000",
x"00000000000000000381f8383f007e03e007c00fc07f03f000060000001fc1f800000000000000003fc003fc0000383c00000000006003f0000000000000",
x"000000000000000003c1f8783f007e03f81f801fc03f83f000040000000fe1f800000000000000003fc003fc00003c380000000001e003f0000000000000",
x"000000000000000003fffff87f80ff033ffe001fc01ffff8000000000007fff800000000000000007f8003fc00001c700000000003e007f0000000000000",
x"000000000000000003fffff9fff7ffc207f8007ff003fffe000000000001ffff0000000000000003ff8001ff800007c0000000000ff81ffe000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007800000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fc00000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013c00000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013c00000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000023800000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040000000000000000000000000",
x"0000000000000000000000000fff8000fff87ffffc7ffffe000f00f07801ffff0001f00010003f03fff0607f83c07ffc004000f81fff1ffe000000000000",
x"00000000000000000000000001fc00001fc0ffffe07ffff8001f83fbfc07fff80007fc003800f3c07f80601e07e00fe000e003fe07fc07f0000000000000",
x"00000000000000000000000001fc00001fc0f80fe07c07f00027c0fcfc1fe1f8000c7e003801e1e03f00700c07e007c000e0063f03fc03f0000000000000",
x"00000000000000000000000000fc00000fc0e007e07003f00007c0f87c3f81f800003f007c03e1e03f00f00c07e007c001f0001f81fc03f0000000000000",
x"00000000000000000000000000fc00000fc0c007e06003f00007c0f87c3f01f800101f007c03e1f03f00f80c03c007c001f0080f80fe03f0000000000000",
x"00000000000000000000000000fc00000fc08007e06003f00007c0f87c7f01f800001f007c03e1f03f01f80c000007c001f8000f807f03f0000000000000",
x"00000000000000000000000000fc00040fc08107e0c003f00007c0f8787f01f800001f80fe07e1f83f01fc0c000007c003f8000fc07f83f0000000000000",
x"00000000000000000000000000fc00040fc08107e0c003f00007c0f8e07f01f800000f80be07c1f83f03fc0c000007c002fc0007c03f83f0000000000000",
x"00000000000000000000000000fc00040fc00107e08003f00007c0f9c07f01f800000f813f07c1f83f03fe0c000007c006fc0007c01fc3f0000000000000",
x"00000000000000000000000000fc00040fc00107e00003f00007c0ff003f01f8001fff813f07c1f83f02fe0c000007c0047c0fffc00fe3f0000000000000",
x"00000000000000000000000000fc00060fc00187e00003f00007c0f8781f81f8001e0f831f87c1f83f067f0c000007c0047e0f07c007f3f0000000000000",
x"00000000000000000000000000fc00078fc001c7e00003f00007c0f87c0fe1f8001e0f021f83e1f03f047f0c000007c0083e0f078007fff0000000000000",
x"00000000000000000000000000fc0007ffc001ffe00003f00007c0f87c07fff8001e0f060f83e1f03f0c3f0c03c007c0083f0f078003fff0000000000000",
x"00000000000000000000000000fc0007ffc001ffe00003f00007c0f87c01fff8000e1e040fc3e1e03f083f8c07e007c0181f070f0001fff0000000000000",
x"00000000000000000000000000fc00070fc001c7e00003f00007c0f83807e1f8000f1e0c07c1e1e03f181f8c07e007c0181f878f0000f3f0000000000000",
x"00000000000000000000000000fc00060fc00187e00003f0007ff87c700fc1f800073c0c0fe0f3c03f181fcc07e007c0381fc39e0000e3f0000000000000",
x"00000000000000000000000000fc00040fc00107e00003f0007fe01fc01f81f80001f01f1ff03f003f301fcc03c007c07e3fe0f8000183f0000000000000",
x"00000000000000000000000000fc00840fc04107e00003f00007c000003f81f800000000000000003f300fec000007c000000000000303f0000000000000",
x"00000000000000000000000100fc04840fc06107e00003f000078000003f81f800000000000000003f200fec000007c000000000000603f0000000000000",
x"00000000000000000000000100fc04840fc06107e00003f000070000003f81f800000000000000003f6007fc000007c000000000001c03f0000000000000",
x"00000000000000000000000180fc0cc00fc06007e00003f000060000001f81f800000000000000003fe007fc000007e400000000003803f0000000000000",
x"000000000000000000000001c0fc1ce00fc07007e00003f000060000001fc1f800000000000000003fc003fc000007f800000000006003f0000000000000",
x"000000000000000000000001e0fc3cf80fc07c07e00003f000040000000fe1f800000000000000003fc003fc000007e00000000001e003f0000000000000",
x"000000000000000000000001fffffcffffc07fffe00007f8000000000007fff800000000000000007f8003fc000007800000000003e007f0000000000000",
x"000000000000000000000001fffffcfffff87ffffc003ffe000000000001ffff0000000000000003ff8001ff80000600000000000ff81ffe000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000780000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000fc0000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000000000000000000013c0000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000000000000000000013c0000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000002380000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000006000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000000000000000",
x"0000000000000000000000000007ffc01fffff00fc107ffffffe0fff80007e00f000001fc004000f81fff1ffe0007cc1f303e001ff003ffe000000000000",
x"0000000000000000000000000000fe003ffff803ff10ffffe0ff01fe0001e781f800007ff00e003fe07fc07f0000e3c38f0ff800fc0007f8000000000000",
x"0000000000000000000000000000fe003e03f80783f0f80fe07f00fc0003c3c27c0001fff00e0063f03fc03f0001c1c70718fc007c0003f0000000000000",
x"00000000000000000000000000007e003801f80f00f0e007e03f80fc0007c3c07c0003c3f01f0001f81fc03f0003c0cf03007e007c0003f0000000000000",
x"00000000000000000000000000007e003001f81e0070c007e01fc0fc0007c3e07c000381f01f0080f80fe03f0003e04f81203e007c0003f0000000000000",
x"00000000000000000000000000007e002001f81e00308007e00fc0fc0007c3e07c000780701f8000f807f03f0003f00fc0003e007c0003f0000000000000",
x"00000000000000000000000000007e002041f81e00108107e00fe0fc000fc3f07c000700003f8000fc07f83f0003fc0ff0003f007c0003f0000000000000",
x"00000000000000000000000000007e002041f81f00108107e007f0fc000f83f07c000f80002fc0007c03f83f0001fe07f8001f007c0003f0000000000000",
x"00000000000000000000000000007e000041f81f80100107e003f8fc000f83f07c000f80006fc0007c01fc3f0001ff07fc001f007c0003f0000000000000",
x"00000000000000000000000000007e000041f81fe0000107e003f8fc000f83f07c000f800047c0fffc00fe3f0000ff83fe3fff007c0003f0000000000000",
x"00000000000000000000000000007e000061f81ff8000187e001fcfc000f83f07c000fc00047e0f07c007f3f00003f80fe3c1f007c0003f0000000000000",
x"00000000000000000000000000007e000071f80ffe0001c7e000fffc0007c3e07c000ff00083e0f078007fff00001fc07f3c1e00fc00fff0000000000000",
x"00000000000000000000000000007e00007ff807ff8001ffe003fffc0007c3e07c0007fc0083f0f078003fff000107c41f3c1e30fc07fff0000000000000",
x"00000000000000000000000000007e00007ff803ffc001ffe00fe0fc0007c3c07c0003ff0181f070f0001fff000183860e1c3c78fc0fe3f0000000000000",
x"00000000000000000000000000007e000071f800ffe001c7e00fc0fc0003c3c07c0001fc0181f878f0000f3f0001c3870e1e3c7d7c1f83f0000000000000",
x"00000000000000000000000000007e000061f8003fe00187e01f80fc0001e787ff8000f00381fc39e0000e3f0001e3078c0e787e7c1f83f0000000000000",
x"00000000000000000000000000007e000041f80007f00107e01f80fc00007e07fe0001e007e3fe0f8000183f00013e04f803e03c7f3f03f0000000000000",
x"00000000000000000000000000007e001041f80803f04107e03f00fc000000007c0003e0000000000000303f0000000000000000003f03f0000000000000",
x"00000000000000000000000000807e021841f80801f06107e03f80fc00000000780003e0000000000000603f0000000000000000003f03f0000000000000",
x"00000000000000000000000000807e021841f80c00f06107e01f80fc00000000700003e0000000000001c03f0000000000000000003f03f0000000000000",
x"00000000000000000000000000c07e061801f80c00f06007e01f80fc00000000600007e0200000000003803f0000000000000000003f83f0000000000000",
x"00000000000000000000000000e07e0e1c01f80f00e07007e01fc0fc00000000600003f0600000000006003f0000000000000000001f83f0000000000000",
x"00000000000000000000000000f07e1e1f01f80f83c07c07e00fe0fc00000000400003ffc0000000001e003f0000000000000000000fe3f0000000000000",
x"00000000000000000000000000fffffe1ffff809ff807fffe007fffe00000000000001ff80000000003e007f00000000000000000007fff8000000000000",
x"00000000000000000000000000fffffe1fffff087e007ffffc00ffff800000000000007e0000000000ff81ffe0000000000000000001fffe000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000780000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000fc0000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000000000000000000013c0000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000000000000000000013c0000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000002380000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000006000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000004000000000000000000000000000000000000000000000000",
x"000000000000000000000000001fff03fc1fff7ffc1ff03ffe000fc100007e00f00007fff004000f81fff1ffe0007cc1f303e001ff003ffe000000000000",
x"0000000000000000000000000003f801fe03fc1fe003c007f0003ff10001e781f80007ffe00e003fe07fc07f0000e3c38f0ff800fc0007f8000000000000",
x"0000000000000000000000000003f800fe01f80fe0018007f000783f0003c3c27c0007ffc00e0063f03fc03f0001c1c70718fc007c0003f0000000000000",
x"0000000000000000000000000001f8007f01f807e0010003f000f00f0007c3c07c0007ffc01f0001f81fc03f0003c0cf03007e007c0003f0000000000000",
x"0000000000000000000000000001f8003f81f807f0030003f001e0070007c3e07c000fff801f0080f80fe03f0003e04f81203e007c0003f0000000000000",
x"0000000000000000000000000001f8001f81f807f0020003f001e0030007c3e07c000c03001f8000f807f03f0003f00fc0003e007c0003f0000000000000",
x"0000000000000000000000000001f8001fc1f803f0060003f001e001000fc3f07c000806003f8000fc07f83f0003fc0ff0003f007c0003f0000000000000",
x"0000000000000000000000000001f8000fe1f803fffe0003f001f001000f83f07c00000c002fc0007c03f83f0001fe07f8001f007c0003f0000000000000",
x"0000000000000000000000000001f80007f1f801fffc0003f001f801000f83f07c00001c006fc0007c01fc3f0001ff07fc001f007c0003f0000000000000",
x"0000000000000000000000000001f80007f1f801fc0c0003f001fe00000f83f07c0000380047c0fffc00fe3f0000ff83fe3fff007c0003f0000000000000",
x"0000000000000000000000000001f80003f9f800fc080003f001ff80000f83f07c0000700047e0f07c007f3f00003f80fe3c1f007c0003f0000000000000",
x"0000000000000000000000000001f80001fff800fc180003f000ffe00007c3e07c0000f00083e0f078007fff00001fc07f3c1e00fc00fff0000000000000",
x"0000000000000000000000000001f80007fff800fe100003f0007ff80007c3e07c0000e00083f0f078003fff000107c41f3c1e30fc07fff0000000000000",
x"0000000000000000000000000001f8001fc1f8007e300003f0003ffc0007c3c07c0001e00181f070f0001fff000183860e1c3c78fc0fe3f0000000000000",
x"0000000000000000000000000001f8001f81f8007f300003f0000ffe0003c3c07c0003e00181f878f0000f3f0001c3870e1e3c7d7c1f83f0000000000000",
x"0000000000000000000000000001f8003f01f8003f600003f00003fe0001e787ff8003e00381fc39e0000e3f0001e3078c0e787e7c1f83f0000000000000",
x"0000000000000000000000000001f8003f01f8003fe00003f000007f00007e07fe0003c007e3fe0f8000183f00013e04f803e03c7f3f03f0000000000000",
x"0000000000000000000000000001f8007e01f8001fc00003f000803f000000007c0007e0000000000000303f0000000000000000003f03f0000000000000",
x"0000000000000000000000000201f8087f01f8001fc00403f010801f00000000780007e0100000000000603f0000000000000000003f03f0000000000000",
x"0000000000000000000000000201f8083f01f8001f800403f010c00f00000000700007e0200000000001c03f0000000000000000003f03f0000000000000",
x"0000000000000000000000000301f8183f01f8000f800603f030c00f00000000600007f8600000000003803f0000000000000000003f83f0000000000000",
x"0000000000000000000000000381f8383f81f8000f800703f070f00e00000000600003ffc00000000006003f0000000000000000001f83f0000000000000",
x"00000000000000000000000003c1f8781fc1f80007000783f0f0f83c00000000400003ffc0000000001e003f0000000000000000000fe3f0000000000000",
x"00000000000000000000000003fffff80ffffc00070007fffff09ff800000000000001ff80000000003e007f00000000000000000007fff8000000000000",
x"00000000000000000000000003fffff801ffff00020007fffff087e0000000000000007e0000000000ff81ffe0000000000000000001fffe000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000001e000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000003f000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000004f000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000004f000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000008e000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000080000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000180000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000001e0f0010003e03fdff7fbffe0ff8001f00fe0001ff7fc1f37fc07fcfe7e01e0f000ff800000000000000000000000",
x"00000000000000000000000000000007f7f803800ff81f8fc3f0ff001e0003fc3ff80007c3f038f1f803f03fff07f7f807fff00000000000000000000000",
x"00000000000000000000000000000001f9f8038018fc1f87c3e07f000c0007fefffc0007c1f07071f001f03f9f01f9f81f81f80000000000000000000000",
x"00000000000000000000000000000001f0f807c0007e1f87c3e03f00080007ffc3fe0007c1f0f031f001f03f0f81f0f83f007e0000000000000000000000",
x"00000000000000000000000000000001f0f807c0203e1f87c3e03f80180008ff80fe0007c1f0f811f001f03e0f81f0f83f003f0000000000000000000000",
x"00000000000000000000000000000001f0f807e0003e1f87c3e03f801000083fc07f0007c1f0fc01f001f03e0f81f0f83f003f8000000000000000000000",
x"00000000000000000000000000000001f0f00fe0003f1f87c3e01f803000001fe07f0007c1f0ff01f001f03e0f81f0f03f001f8000000000000000000000",
x"00000000000000000000000000000001f1c00bf0001f1f87c3e01ffff000003ff03e0007c1f07f81f001f03e0f81f1c03f001fc000000000000000000000",
x"00000000000000000000000000000001f3801bf0001f1f87c3e00fffe0000067f03e0007c1f07fc1f001f03e0f81f3803f000fc000000000000000000000",
x"00000000000000000000000000000001fe0011f03fff1f87c3e00fe060000063f83e0007c1f03fe1f001f03e0f81fe007f800fc000000000000000000000",
x"00000000000000000000000000000001f0f011f83c1f1f87c3e007e0400000c1fc3c0007c1f00fe1f001f03e0f81f0f1ffe00fc000000000000000000000",
x"00000000000000000000000000000001f0f820f83c1e1f87c3e007e0c00001c0fc380007c1f007f1f003f03e0f81f0f800000fe000000000000000000000",
x"00000000000000000000000000000001f0f820fc3c1e1f87c3e007f0800001c0fee00007c1f041f1f0c3f03e0f81f0f800000fe000000000000000000000",
x"00000000000000000000000000000001f0f8607c1c3c1f8fc3e003f1800003c07f800007c3f060e1f1e3f03e0f81f0f800000fc000000000000000000000",
x"00000000000000000000000000000001f070607e1e3c0f9fe7e003f980000ff03f000007e7f070e1f1f5f03e0f81f07000000fc000000000000000000000",
x"00000000000000000000000000000000f8e0e07f0e780ff3fbf001fb000000007f000003fdf078c1f9f9f03f0f80f8e000000fc000000000000000000000",
x"000000000000000000000000000000003f81f8ff83e007c1f3f801ff00000001df000001f1f04f81fcf1fc3f8fe03f8000001fc000000000000000000000",
x"000000000000000000000000000000000000000000000000000000fe000000071f80000001f00000000000000000000020001f8000000000000000000000",
x"000000000000000000000000000000000000000000000000000000fe0000000f0f80000001f00000000000000000000030001f8000000000000000000000",
x"000000000000000000000000000000000000000000000000000000fc0000000f0f80000001f00000000000000000000030003f0000000000000000000000",
x"0000000000000000000000000000000000000000000000000000007c0000000f0f00000001f00000e00000000000000038003e0000000000000000000000",
x"0000000000000000000000000000000000000000000000000000007c0000000f0f00000001f00001f0000000000000003e007c0000000000000000000000",
x"000000000000000000000000000000000000000000000000000000380000000f0e00000001f00001f8000000000000003f81f80000000000000000000000",
x"00000000000000000000000000000000000000000000000000000038000000078c00000001f00001f00000000000000033ffe00000000000000000000000",
x"0000000000000000000000000000000000000000000000000000001000000003f000000001fc0000e000000000000000207f800000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000007ffe000ffff80000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000fe0003fffc00000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000fe000ff0fc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000007e001fc0fc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000007e001f80fc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000007e003f80fc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000007e003f80fc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000007e003f80fc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000007e003f80fc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000007e001f80fc00000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000fe000fc0fc00000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000ff0007f0fc00000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000001bf0003fffc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000013f8000fffc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000031f8003f0fc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000061fc007e0fc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000060fc00fc0fc00000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000c07e01fc0fc00000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000807f01fc0fc00000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000001803f01fc0fc00000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000003003f80fc0fc00000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000003001f80fe0fc00000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000007001fc07f0fc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000000f001fe03fffc00000000000000000000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000000000000000000001fc07ff80ffff80000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000ff81f03f9ff0f07807c003fe01ffff003f9ff03e07fc07fc03fffe000000000000000000000000000000000000",
x"00000000000000000000000000000000007e07fc1f8fe3fbfc1ff001f807fff8001f8fe0ff81f803f00ffff0000000000000000000000000000000000000",
x"00000000000000000000000000000000003e0c7e0f87c0fcfc31f800f81fe1f8000f87c10fc1f001f03fc3f0000000000000000000000000000000000000",
x"00000000000000000000000000000000003e003f0f87c0f87c00fc00f83f81f8000f87c207e1f001f07f03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000003e101f07c7c0f87c407c00f83f01f80007c7c007e1f001f07e03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000003e001f07e7c0f87c007c00f87f01f80007e7c003e1f001f0fe03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000003e001f83e7c0f878007e00f87f01f80003e7c003f1f001f0fe03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000003e000f81ffc0f8e0003e00f87f01f80001ffc003f1f001f0fe03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000003e000f81ffc0f9c0003e00f87f01f80001ffc001f1f001f0fe03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000003e1fff80f7c0ff007ffe00f83f01f80000f7c001f1f001f07e03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000003e1e0f8067c0f878783e00f81f81f8000067c001f1f001f03f03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000007e1e0f0047c0f87c783c01f80fe1f8000047c001e1f003f01fc3f0000000000000000000000000000000000000",
x"00000000000000000000000000000000187e1e0f0087c0f87c783c61f807fff8000087c1c1e1f0c3f00ffff0000000000000000000000000000000000000",
x"000000000000000000000000000000003c7e0e1e0107c0f87c3878f1f801fff8000107c3e3c1f1e3f003fff0000000000000000000000000000000000000",
x"000000000000000000000000000000003ebe0f1e0307c0f8383c78faf807e1f8000307c3e3c1f1f5f00fc3f0000000000000000000000000000000000000",
x"000000000000000000000000000000003f3e073c0707c07c701cf0fcf80fc1f8000707c1e781f9f9f01f83f0000000000000000000000000000000000000",
x"000000000000000000000000000000001e3f81f01fc7c01fc007c078fe1f81f8001fc7c07e01fcf1fc3f03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000007c00000000000003f81f8000007c000000000007f03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000007c00000000000003f81f8000007c000000000007f03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000007c00000000000003f81f8000007c000000000007f03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000007c00000000000001f81f8000007c00000e000003f03f0000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000007c00000000000001fc1f8000007c00001f000003f83f0000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000007c00000000000000fe1f8000007c00001f800001fc3f0000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000007e000000000000007fff8000007e00001f000000ffff0000000000000000000000000000000000000",
x"00000000000000000000000000000000000000000007f000000000000001ffff000007f00000e0000003fffe000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
);
	
	

constant paused_rom: rom_paused :=
	(
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000003ff8000c00000001fff800000000000000000000000000000000000000",
x"00000000fffffffff807fffffffffffff00001ffff000c0000001fffff8000007fffffff0001fffff0000007fffffffc",
x"0000001ffffffffff807fffffffffffff00007ffffe01c0000007fffffe000007fffffff0001fffff0000007fffffffc",
x"000000fffffffffe0007fffffffffffe00001ff00ff87c000001fffffff800001fffffc000001fffc00000003fffff00",
x"000003ffe03ffffc0007fff0007ffff800007fc001fffc000003f803fffc000007ffff80000003ff000000000ffffc00",
x"00000fff000ffff8000fff80003ffff00000ff00007ffc000007c000ffff000003ffff00000001fe0000000007fffc00",
x"00003ffe000ffff0000ffe00001fffe00001fe00003ffc00001f80003fff800001ffff00000001fc0000000007fff800",
x"00007ff8000ffff0000ff800001fffe00003fc00000ffc00001e00001fff800000ffff00000001f80000000003fff800",
x"0001fff0000ffff0000ff000001fffe00007fc000007fc00003c00000fffc00000ffff80000001f80000000003fff800",
x"0003fff0000ffff0000fe000000fffe00007f8000003fc00007800000fffe000007fff80000001f00000000003fff800",
x"0007ffe0000ffff0000fc000000fffe0000ff8000001fc0000f8000007ffe000007fffc0000001f00000000003fff800",
x"000fffc0000ffff0000f8000000fffe0000ff8000001fc0000f0000007fff000003fffc0000001e00000000003fff800",
x"001fffc0000ffff0001f0000000fffe0001ff8000000fc0001f0000007fff000003fffc0000003e00000000003fff800",
x"001fff80000ffff0001e0000000fffe0001ff80000007c0001e0000003fff800001fffe0000003c00000000003fff800",
x"003fff80000ffff0001e0000000fffe0001ff80000007c0001e0000003fff800001fffe0000007c00000000003fff800",
x"007fff80000ffff0001c0000000fffe0003ff80000003c0001e0000003fff800000ffff0000007800000000003fff800",
x"007fff00000ffff0001c0000000fffe0003ffc0000003c0003c0000003fff800000ffff0000007800000000003fff800",
x"00ffff00000ffff00018000c000fffe0003ffc0000001c0003c0000003fff800000ffff800000f000000000003fff800",
x"00ffff00000ffff00018000c000fffe0003ffe0000001c0003c0000003fff8000007fff800000f000000000003fff800",
x"01fffe00000ffff00038000e000fffe0003fff0000001c0003c0000003fffc000007fffffffffe000000000003fff800",
x"01fffe00000ffff00030000e000fffe0003fff8000000c0003c0000003fffc000003fffffffffe000000000003fff800",
x"01fffe00000ffff00000000e000fffe0003fffc000000c0003c0000003fffc000003fffffffffc000000000003fff800",
x"03fffe00000ffff00000000e000fffe0003ffff000000c0003c0000003fffc000001fffffffffc000000000003fff800",
x"03fffe00000ffff00000000f000fffe0003ffff800000c0003c0000003fffc000001fffe00007c000000000003fff800",
x"03fffe00000ffff00000000f000fffe0001ffffe0000000003c0000003fffc000001ffff000078000000000003fff800",
x"03fffc00000ffff00000000f000fffe0001fffff8000000003c0000003fffc000000ffff000078000000000003fff800",
x"07fffc00000ffff00000000f800fffe0001fffffe000000003c0000003fffc000000ffff0000f0000000000003fff800",
x"07fffc00000ffff00000000f800fffe0000ffffff800000003c0000003fffc0000007fff8000f0000000000003fff800",
x"07fffc00000ffff00000000fc00fffe0000ffffffe00000003c0000003fffc0000007fff8001e0000000000003fff800",
x"07fffc00000ffff00000000fe00fffe00007ffffff80000003c0000003fffc0000003fffc001e0000000000003fff800",
x"07fffc00000ffff00000000ff00fffe00003ffffffc0000003c0000003fffc0000003fffc003c0000000000003fff800",
x"07fffc00000ffff00000000ffe0fffe00001fffffff0000003c0000003fffc0000001fffe003c0000000003ffffff800",
x"07fffc00000ffff00000000fffffffe00000fffffff8000003c0000003fffc0000001fffe007c000000007fffffff800",
x"07fffc00000ffff00000000fffffffe000007ffffffe000003c0000003fffc0000001fffe007800000003ffffffff800",
x"07fffc00000ffff00000000fffffffe000003fffffff000003c0000003fffc0000000ffff00f80000000fffe03fff800",
x"07fffc00000ffff00000000ffe0fffe000001fffffff800003c0000003fffc0000000ffff00f00000001fff803fff800",
x"07fffc00000ffff00000000ff00fffe0000007ffffffc00003c0000003fffc00000007fff80f00000007fff003fff800",
x"07fffc00000ffff00000000fe00fffe0000001ffffffe00003c0000003fffc00000007fff81e0000000fffe003fff800",
x"07fffc00000ffff00000000fc00fffe0000000ffffffe00003c0000003fffc00000003fffc1e0000001fffc003fff800",
x"07fffc00000ffff00000000f800fffe00000003ffffff00003c0000003fffc00000003fffc3c0000001fff8003fff800",
x"03fffe00000ffff00000000f800fffe00000000ffffff00003c0000003fffc00000003fffc3c0000003fff8003fff800",
x"03fffe00000ffff00000000f000fffe000000003fffff80003c0000003fffc00000001fffe7c0000007fff8003fff800",
x"03fffe00000ffff00000000f000fffe000000000fffff80003c0000003fffc00000001fffe780000007fff0003fff800",
x"03fffe00000ffff00000000f000fffe0000000003ffffc0003c0000003fffc00000000fffff80000007fff0003fff800",
x"01fffe00000ffff00000000e000fffe0000000000ffffc0003c0000003fffc00000000fffff0000000ffff0003fff800",
x"01fffe00000ffff00000000e000fffe00003000007fffc0003c0000003fffc000000007ffff0000000ffff0003fff800",
x"01ffff00000ffff00001800e000fffe00003000001fffc0003c0000003fffc000000007fffe0000000ffff0003fff800",
x"00ffff00000ffff00001800e000fffe00003000000fffc0003c0000003fffc000000007fffe0000000ffff0003fff800",
x"00ffff00000ffff00001800c000fffe000038000007ffc0003c0000003fffc000000003fffc0000000ffff0003fff800",
x"007fff80000ffff00001800c000fffe000038000003ffc0003c0000003fffc000000003fffc0000000ffff0003fff800",
x"007fff80000ffff00001c000000fffe000038000001ffc0003c0000003fffc000000001fffc0000000ffff0003fff800",
x"003fff80000ffff00001c000000fffe00003c000001ffc0003c0000003fffc000000001fff80000000ffff0003fff800",
x"001fffc0000ffff00001e000000fffe00003c000000ffc0003c0000003fffc000000000fff80000000ffff0003fff800",
x"001fffc0000ffff00001e000000fffe00003e000000ff80003c0000003fffc000000000fff000000007fff0003fff800",
x"000fffe0000ffff00001f000000fffe00003e000000ff80003c0000003fffc000000000fff000000007fff0003fff800",
x"0007fff0000ffff00001f000000fffe00003f000000ff00003c0000003fffc0000000007fe000000003fff8003fff800",
x"0003fff0000ffff00001f800000fffe00003f800000ff00007c0000003fffc0000000007fe000000003fff8003fff800",
x"0001fff8000ffff00001fc00000fffe00003fc00001fe00007c0000003fffc0000000003fc000000001fffc003fff800",
x"0000fffc000ffff00001ff00000fffe00003fe00001fe00007c0000003fffc0000000003fc000000000fffe003fff800",
x"00003fff000ffff00001ffc0000fffe00003ff00003fc00007c0000003fffc0000000001fc0000000007fff003fff800",
x"00001fff800ffff80001fff8000ffff00003ffc0007f80000fe0000003fffc0000000001f80000000003fff803fffc00",
x"000007fff80ffffc0001fffffffffff80003ffe000ff00001ff0000007fffe0000000000f80000000000ffff03fffc00",
x"000000fffffffffe0001fffffffffffe000387fc07fe00007ffc00001fffff8000000000f000000000003fffffffff00",
x"0000001ffffffffff801fffffffffffff00380fffff80007ffffe007fffffffc00000000f0000000000007fffffffffc",
x"00000000fffffffff801fffffffffffff003003fffe00007ffffe007fffffffc00000000600000000000003ffffffffc",
x"0000000000000000000000000000000000030007ff000000000000000000000000000000600000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
x"000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
);

constant ball_rom: rom_ball :=
	(
		"0000000000000",
		"0000000000000",
		"0000000000000",
		"0000111110000",
		"0001111111000",
		"0011111111100",
		"0011111111100",
		"0011111111100",
		"0011111111100",
		"0001111111000",
		"0000111110000",
		"0000000000000",
		"0000000000000"
);

	begin
		
		ball_single_row <= ball_rom(ball_row);--to determine which pixel to color with ball color
		ball_validity_bit <= ball_single_row(ball_col);
					
		r_ball<="0000";--ball color
		g_ball<="1111";
		b_ball<="0000";
		
		welmes_single_row <= welmes_rom(welmes_row);--to determine which pixel to color with welcome message color
		welmes_validity_bit <= welmes_single_row(welmes_col);
					
		r_welmes<="1111";--welcome message color
		g_welmes<="1111";
		b_welmes<="0000";
		
		paused_single_row <= paused_rom(paused_row);--to determine which pixel to color with pause message color
		paused_validity_bit <= paused_single_row(paused_col);
					
		r_paused<="1111";--pause message color
		g_paused<="1000";
		b_paused<="0000";
		
		winmes_single_row <= winmes_rom(winmes_row);--to determine which pixel to color with win message color
		winmes_validity_bit <= winmes_single_row(winmes_col);
					
		r_winmes<="0000";--win message color
		g_winmes<="0000";
		b_winmes<="1111";
		
		gameover_single_row <= gameover_rom(gameover_row);--to determine which pixel to color with gameover message color
		gameover_validity_bit <= gameover_single_row(gameover_col);
					
		r_gameover<="1111";--gameover message color
		g_gameover<="0000";
		b_gameover<="0000";
		
		lives_single_row <=lives3_rom(lives_row)when isalive=3 else--to determine which pixel to color with lives message color
								 lives2_rom(lives_row)when isalive=2 else
								 lives1_rom(lives_row)when isalive=1 else
							    lives0_rom(lives_row);
		
		lives_validity_bit <= lives_single_row(lives_col);
					
		r_lives<="0000";--lives message color
		g_lives<="1111";
		b_lives<="1111";
		
		hpos_scr<=hpos-152 when (hpos>152 and hpos<793)else
					 1;--bring x and y position inside screen by
		vpos_scr<=vpos-37 when (vpos>37 and vpos<518)else
					 1;--subtracting fp,bp and sync period
		
		process(clk_s)--process to generate random postion of x for ball and bat
			begin
				
				if(clk_s'event and clk_s='0') then
					ball_x_vel_rand<=not ball_x_vel_rand;
					if(rand_x=611)then
						rand_x<=26;
					else
						rand_x<=rand_x+3;
					end if;
				end if;
		end process;
		
		process(clk_s)--main synchronization process
			begin
				
				if(clk_s'event and clk_s='1') then									
														
					if(resetgame='0') then--to reset game after key3 has been pressed
						notstarted<='1';
						isalive<=3;
						ball_x<=rand_x;
						ball_y<=450;
						bat_x<=rand_x-25;
						bat_y<=460;
						ball_x_vel<=ball_x_vel_rand;
						ball_y_vel<='0';
						is_destroyed_l1<=x"000000000000000000";
						coll_x_l1<=x"000000000000000000";
						coll_y_l1<=x"000000000000000000";
						is_destroyed_l2<=x"0000000";
						coll_x_l2<=x"0000000";
						coll_y_l2<=x"0000000";
						is_destroyed_l3<=x"000000000000000000";
						coll_x_l3<=x"000000000000000000";
						coll_y_l3<=x"000000000000000000";
						is_destroyed_l4<=x"0000000000000000";
						coll_x_l4<=x"0000000000000000";
						coll_y_l4<=x"0000000000000000";
						is_destroyed_l5<=x"000000000";
						coll_x_l5<=x"000000000";
						coll_y_l5<=x"000000000";
						l1complete<='0';
						l2complete<='0';
						l3complete<='0';
						l4complete<='0';
						l5complete<='0';
						l2notstarted<='1';
						l3notstarted<='1';
						l4notstarted<='1';
						l5notstarted<='1';
						level_selected<='0';
						stopball<='0';
					else
						null;
					end if;
					
					if(level_selected='0')then--to select level at the start of the game
						case level_select is
							when "010"=>l1complete<='1';
											l2complete<='0';
											l3complete<='0';
											l4complete<='0';
											l5complete<='0';
											l2notstarted<='0';
											l3notstarted<='1';
											l4notstarted<='1';
											l5notstarted<='1';
							when "011"=>l1complete<='1';
											l2complete<='1';
											l3complete<='0';
											l4complete<='0';
											l5complete<='0';
											l2notstarted<='0';
											l3notstarted<='0';
											l4notstarted<='1';
											l5notstarted<='1';
							when "100"=>l1complete<='1';
											l2complete<='1';
											l3complete<='1';
											l4complete<='0';
											l5complete<='0';
											l2notstarted<='0';
											l3notstarted<='0';
											l4notstarted<='0';
											l5notstarted<='1';
							when "101"=>l1complete<='1';
											l2complete<='1';
											l3complete<='1';
											l4complete<='1';
											l5complete<='0';
											l2notstarted<='0';
											l3notstarted<='0';
											l4notstarted<='0';
											l5notstarted<='0';
							when others=>l1complete<='0';
											l2complete<='0';
											l3complete<='0';
											l4complete<='0';
											l5complete<='0';
											l2notstarted<='1';
											l3notstarted<='1';
											l4notstarted<='1';
											l5notstarted<='1';
						end case;
					else
						null;
					end if;
					
					
					if(l2notstarted='1'and is_destroyed_l1=x"ffffffffffffffffff")then--to start level 2
						ball_x<=rand_x;
						ball_y<=450;
						bat_x<=rand_x-25;
						bat_y<=460;
						ball_x_vel<=ball_x_vel_rand;
						ball_y_vel<='0';
						l1complete<='1';
						l2notstarted<='0';
					elsif(l3notstarted='1'and is_destroyed_l2=x"fffffff")then--to start level 3
						ball_x<=rand_x;
						ball_y<=450;
						bat_x<=rand_x-25;
						bat_y<=460;
						ball_x_vel<=ball_x_vel_rand;
						ball_y_vel<='0';
						l2complete<='1';
						l3notstarted<='0';
					elsif(l4notstarted='1'and is_destroyed_l3=x"ffffffffffffffffff")then--to start level 4
						ball_x<=rand_x;
						ball_y<=450;
						bat_x<=rand_x-25;
						bat_y<=460;
						ball_x_vel<=ball_x_vel_rand;
						ball_y_vel<='0';
						l3complete<='1';
						l4notstarted<='0';
					elsif(l5notstarted='1'and is_destroyed_l4=x"ffffffffffffffff")then--to start level 5
						ball_x<=rand_x;
						ball_y<=450;
						bat_x<=rand_x-25;
						bat_y<=460;
						ball_x_vel<=ball_x_vel_rand;
						ball_y_vel<='0';
						l4complete<='1';
						l5notstarted<='0';
					elsif(is_destroyed_l5=x"fffffffff")then--to complete level 5
						l5complete<='1';
					else 
						null;
					end if;

					if(start='0' and level_select/="000" and level_select/="110" and level_select/="111") then--start the game and stop level selection only if valid level is selected
						notstarted<='0';
						level_selected<='1';
					else
						null;
					end if;
					
					if(notstarted='0') then
						if(l1complete='0')then--display bricks of level 1
							brick(hpos_scr,vpos_scr,x_cood_l1(71),y_cood_l1(71),ball_x,ball_y,draw_l1(71),r_brick(71),g_brick(71),b_brick(71),coll_x_l1(71),coll_y_l1(71),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(70),y_cood_l1(70),ball_x,ball_y,draw_l1(70),r_brick(70),g_brick(70),b_brick(70),coll_x_l1(70),coll_y_l1(70),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(69),y_cood_l1(69),ball_x,ball_y,draw_l1(69),r_brick(69),g_brick(69),b_brick(69),coll_x_l1(69),coll_y_l1(69),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(68),y_cood_l1(68),ball_x,ball_y,draw_l1(68),r_brick(68),g_brick(68),b_brick(68),coll_x_l1(68),coll_y_l1(68),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(67),y_cood_l1(67),ball_x,ball_y,draw_l1(67),r_brick(67),g_brick(67),b_brick(67),coll_x_l1(67),coll_y_l1(67),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(66),y_cood_l1(66),ball_x,ball_y,draw_l1(66),r_brick(66),g_brick(66),b_brick(66),coll_x_l1(66),coll_y_l1(66),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(65),y_cood_l1(65),ball_x,ball_y,draw_l1(65),r_brick(65),g_brick(65),b_brick(65),coll_x_l1(65),coll_y_l1(65),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(64),y_cood_l1(64),ball_x,ball_y,draw_l1(64),r_brick(64),g_brick(64),b_brick(64),coll_x_l1(64),coll_y_l1(64),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(63),y_cood_l1(63),ball_x,ball_y,draw_l1(63),r_brick(63),g_brick(63),b_brick(63),coll_x_l1(63),coll_y_l1(63),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(62),y_cood_l1(62),ball_x,ball_y,draw_l1(62),r_brick(62),g_brick(62),b_brick(62),coll_x_l1(62),coll_y_l1(62),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(61),y_cood_l1(61),ball_x,ball_y,draw_l1(61),r_brick(61),g_brick(61),b_brick(61),coll_x_l1(61),coll_y_l1(61),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(60),y_cood_l1(60),ball_x,ball_y,draw_l1(60),r_brick(60),g_brick(60),b_brick(60),coll_x_l1(60),coll_y_l1(60),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(59),y_cood_l1(59),ball_x,ball_y,draw_l1(59),r_brick(59),g_brick(59),b_brick(59),coll_x_l1(59),coll_y_l1(59),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(58),y_cood_l1(58),ball_x,ball_y,draw_l1(58),r_brick(58),g_brick(58),b_brick(58),coll_x_l1(58),coll_y_l1(58),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(57),y_cood_l1(57),ball_x,ball_y,draw_l1(57),r_brick(57),g_brick(57),b_brick(57),coll_x_l1(57),coll_y_l1(57),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(56),y_cood_l1(56),ball_x,ball_y,draw_l1(56),r_brick(56),g_brick(56),b_brick(56),coll_x_l1(56),coll_y_l1(56),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(55),y_cood_l1(55),ball_x,ball_y,draw_l1(55),r_brick(55),g_brick(55),b_brick(55),coll_x_l1(55),coll_y_l1(55),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(54),y_cood_l1(54),ball_x,ball_y,draw_l1(54),r_brick(54),g_brick(54),b_brick(54),coll_x_l1(54),coll_y_l1(54),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(53),y_cood_l1(53),ball_x,ball_y,draw_l1(53),r_brick(53),g_brick(53),b_brick(53),coll_x_l1(53),coll_y_l1(53),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(52),y_cood_l1(52),ball_x,ball_y,draw_l1(52),r_brick(52),g_brick(52),b_brick(52),coll_x_l1(52),coll_y_l1(52),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(51),y_cood_l1(51),ball_x,ball_y,draw_l1(51),r_brick(51),g_brick(51),b_brick(51),coll_x_l1(51),coll_y_l1(51),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(50),y_cood_l1(50),ball_x,ball_y,draw_l1(50),r_brick(50),g_brick(50),b_brick(50),coll_x_l1(50),coll_y_l1(50),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(49),y_cood_l1(49),ball_x,ball_y,draw_l1(49),r_brick(49),g_brick(49),b_brick(49),coll_x_l1(49),coll_y_l1(49),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(48),y_cood_l1(48),ball_x,ball_y,draw_l1(48),r_brick(48),g_brick(48),b_brick(48),coll_x_l1(48),coll_y_l1(48),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(47),y_cood_l1(47),ball_x,ball_y,draw_l1(47),r_brick(47),g_brick(47),b_brick(47),coll_x_l1(47),coll_y_l1(47),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(46),y_cood_l1(46),ball_x,ball_y,draw_l1(46),r_brick(46),g_brick(46),b_brick(46),coll_x_l1(46),coll_y_l1(46),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(45),y_cood_l1(45),ball_x,ball_y,draw_l1(45),r_brick(45),g_brick(45),b_brick(45),coll_x_l1(45),coll_y_l1(45),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(44),y_cood_l1(44),ball_x,ball_y,draw_l1(44),r_brick(44),g_brick(44),b_brick(44),coll_x_l1(44),coll_y_l1(44),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(43),y_cood_l1(43),ball_x,ball_y,draw_l1(43),r_brick(43),g_brick(43),b_brick(43),coll_x_l1(43),coll_y_l1(43),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(42),y_cood_l1(42),ball_x,ball_y,draw_l1(42),r_brick(42),g_brick(42),b_brick(42),coll_x_l1(42),coll_y_l1(42),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(41),y_cood_l1(41),ball_x,ball_y,draw_l1(41),r_brick(41),g_brick(41),b_brick(41),coll_x_l1(41),coll_y_l1(41),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(40),y_cood_l1(40),ball_x,ball_y,draw_l1(40),r_brick(40),g_brick(40),b_brick(40),coll_x_l1(40),coll_y_l1(40),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(39),y_cood_l1(39),ball_x,ball_y,draw_l1(39),r_brick(39),g_brick(39),b_brick(39),coll_x_l1(39),coll_y_l1(39),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(38),y_cood_l1(38),ball_x,ball_y,draw_l1(38),r_brick(38),g_brick(38),b_brick(38),coll_x_l1(38),coll_y_l1(38),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(37),y_cood_l1(37),ball_x,ball_y,draw_l1(37),r_brick(37),g_brick(37),b_brick(37),coll_x_l1(37),coll_y_l1(37),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(36),y_cood_l1(36),ball_x,ball_y,draw_l1(36),r_brick(36),g_brick(36),b_brick(36),coll_x_l1(36),coll_y_l1(36),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(35),y_cood_l1(35),ball_x,ball_y,draw_l1(35),r_brick(35),g_brick(35),b_brick(35),coll_x_l1(35),coll_y_l1(35),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(34),y_cood_l1(34),ball_x,ball_y,draw_l1(34),r_brick(34),g_brick(34),b_brick(34),coll_x_l1(34),coll_y_l1(34),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(33),y_cood_l1(33),ball_x,ball_y,draw_l1(33),r_brick(33),g_brick(33),b_brick(33),coll_x_l1(33),coll_y_l1(33),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(32),y_cood_l1(32),ball_x,ball_y,draw_l1(32),r_brick(32),g_brick(32),b_brick(32),coll_x_l1(32),coll_y_l1(32),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(31),y_cood_l1(31),ball_x,ball_y,draw_l1(31),r_brick(31),g_brick(31),b_brick(31),coll_x_l1(31),coll_y_l1(31),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(30),y_cood_l1(30),ball_x,ball_y,draw_l1(30),r_brick(30),g_brick(30),b_brick(30),coll_x_l1(30),coll_y_l1(30),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(29),y_cood_l1(29),ball_x,ball_y,draw_l1(29),r_brick(29),g_brick(29),b_brick(29),coll_x_l1(29),coll_y_l1(29),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(28),y_cood_l1(28),ball_x,ball_y,draw_l1(28),r_brick(28),g_brick(28),b_brick(28),coll_x_l1(28),coll_y_l1(28),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(27),y_cood_l1(27),ball_x,ball_y,draw_l1(27),r_brick(27),g_brick(27),b_brick(27),coll_x_l1(27),coll_y_l1(27),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(26),y_cood_l1(26),ball_x,ball_y,draw_l1(26),r_brick(26),g_brick(26),b_brick(26),coll_x_l1(26),coll_y_l1(26),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(25),y_cood_l1(25),ball_x,ball_y,draw_l1(25),r_brick(25),g_brick(25),b_brick(25),coll_x_l1(25),coll_y_l1(25),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(24),y_cood_l1(24),ball_x,ball_y,draw_l1(24),r_brick(24),g_brick(24),b_brick(24),coll_x_l1(24),coll_y_l1(24),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(23),y_cood_l1(23),ball_x,ball_y,draw_l1(23),r_brick(23),g_brick(23),b_brick(23),coll_x_l1(23),coll_y_l1(23),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(22),y_cood_l1(22),ball_x,ball_y,draw_l1(22),r_brick(22),g_brick(22),b_brick(22),coll_x_l1(22),coll_y_l1(22),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(21),y_cood_l1(21),ball_x,ball_y,draw_l1(21),r_brick(21),g_brick(21),b_brick(21),coll_x_l1(21),coll_y_l1(21),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(20),y_cood_l1(20),ball_x,ball_y,draw_l1(20),r_brick(20),g_brick(20),b_brick(20),coll_x_l1(20),coll_y_l1(20),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(19),y_cood_l1(19),ball_x,ball_y,draw_l1(19),r_brick(19),g_brick(19),b_brick(19),coll_x_l1(19),coll_y_l1(19),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(18),y_cood_l1(18),ball_x,ball_y,draw_l1(18),r_brick(18),g_brick(18),b_brick(18),coll_x_l1(18),coll_y_l1(18),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(17),y_cood_l1(17),ball_x,ball_y,draw_l1(17),r_brick(17),g_brick(17),b_brick(17),coll_x_l1(17),coll_y_l1(17),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(16),y_cood_l1(16),ball_x,ball_y,draw_l1(16),r_brick(16),g_brick(16),b_brick(16),coll_x_l1(16),coll_y_l1(16),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(15),y_cood_l1(15),ball_x,ball_y,draw_l1(15),r_brick(15),g_brick(15),b_brick(15),coll_x_l1(15),coll_y_l1(15),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(14),y_cood_l1(14),ball_x,ball_y,draw_l1(14),r_brick(14),g_brick(14),b_brick(14),coll_x_l1(14),coll_y_l1(14),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(13),y_cood_l1(13),ball_x,ball_y,draw_l1(13),r_brick(13),g_brick(13),b_brick(13),coll_x_l1(13),coll_y_l1(13),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(12),y_cood_l1(12),ball_x,ball_y,draw_l1(12),r_brick(12),g_brick(12),b_brick(12),coll_x_l1(12),coll_y_l1(12),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(11),y_cood_l1(11),ball_x,ball_y,draw_l1(11),r_brick(11),g_brick(11),b_brick(11),coll_x_l1(11),coll_y_l1(11),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(10),y_cood_l1(10),ball_x,ball_y,draw_l1(10),r_brick(10),g_brick(10),b_brick(10),coll_x_l1(10),coll_y_l1(10),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(9),y_cood_l1(9),ball_x,ball_y,draw_l1(9),r_brick(9),g_brick(9),b_brick(9),coll_x_l1(9),coll_y_l1(9),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(8),y_cood_l1(8),ball_x,ball_y,draw_l1(8),r_brick(8),g_brick(8),b_brick(8),coll_x_l1(8),coll_y_l1(8),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(7),y_cood_l1(7),ball_x,ball_y,draw_l1(7),r_brick(7),g_brick(7),b_brick(7),coll_x_l1(7),coll_y_l1(7),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(6),y_cood_l1(6),ball_x,ball_y,draw_l1(6),r_brick(6),g_brick(6),b_brick(6),coll_x_l1(6),coll_y_l1(6),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(5),y_cood_l1(5),ball_x,ball_y,draw_l1(5),r_brick(5),g_brick(5),b_brick(5),coll_x_l1(5),coll_y_l1(5),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(4),y_cood_l1(4),ball_x,ball_y,draw_l1(4),r_brick(4),g_brick(4),b_brick(4),coll_x_l1(4),coll_y_l1(4),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(3),y_cood_l1(3),ball_x,ball_y,draw_l1(3),r_brick(3),g_brick(3),b_brick(3),coll_x_l1(3),coll_y_l1(3),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(2),y_cood_l1(2),ball_x,ball_y,draw_l1(2),r_brick(2),g_brick(2),b_brick(2),coll_x_l1(2),coll_y_l1(2),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(1),y_cood_l1(1),ball_x,ball_y,draw_l1(1),r_brick(1),g_brick(1),b_brick(1),coll_x_l1(1),coll_y_l1(1),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l1(0),y_cood_l1(0),ball_x,ball_y,draw_l1(0),r_brick(0),g_brick(0),b_brick(0),coll_x_l1(0),coll_y_l1(0),ball_x_vel,ball_y_vel);
							ball(hpos_scr,vpos_scr,ball_x,ball_y,ball_row,ball_col);	--get the ball image
						elsif(l2complete='0')then--display bricks of level 2
							brick(hpos_scr,vpos_scr,x_cood_l2(71),y_cood_l2(71),ball_x,ball_y,draw_l2(71),r_brick(71),g_brick(71),b_brick(71),coll_x_l2(71),coll_y_l2(71),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(70),y_cood_l2(70),ball_x,ball_y,draw_l2(70),r_brick(70),g_brick(70),b_brick(70),coll_x_l2(70),coll_y_l2(70),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(69),y_cood_l2(69),ball_x,ball_y,draw_l2(69),r_brick(69),g_brick(69),b_brick(69),coll_x_l2(69),coll_y_l2(69),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(68),y_cood_l2(68),ball_x,ball_y,draw_l2(68),r_brick(68),g_brick(68),b_brick(68),coll_x_l2(68),coll_y_l2(68),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(67),y_cood_l2(67),ball_x,ball_y,draw_l2(67),r_brick(67),g_brick(67),b_brick(67),coll_x_l2(67),coll_y_l2(67),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(66),y_cood_l2(66),ball_x,ball_y,draw_l2(66),r_brick(66),g_brick(66),b_brick(66),coll_x_l2(66),coll_y_l2(66),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(65),y_cood_l2(65),ball_x,ball_y,draw_l2(65),r_brick(65),g_brick(65),b_brick(65),coll_x_l2(65),coll_y_l2(65),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(64),y_cood_l2(64),ball_x,ball_y,draw_l2(64),r_brick(64),g_brick(64),b_brick(64),coll_x_l2(64),coll_y_l2(64),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(63),y_cood_l2(63),ball_x,ball_y,draw_l2(63),r_brick(63),g_brick(63),b_brick(63),coll_x_l2(63),coll_y_l2(63),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(62),y_cood_l2(62),ball_x,ball_y,draw_l2(62),r_brick(62),g_brick(62),b_brick(62),coll_x_l2(62),coll_y_l2(62),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(61),y_cood_l2(61),ball_x,ball_y,draw_l2(61),r_brick(61),g_brick(61),b_brick(61),coll_x_l2(61),coll_y_l2(61),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(60),y_cood_l2(60),ball_x,ball_y,draw_l2(60),r_brick(60),g_brick(60),b_brick(60),coll_x_l2(60),coll_y_l2(60),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(59),y_cood_l2(59),ball_x,ball_y,draw_l2(59),r_brick(59),g_brick(59),b_brick(59),coll_x_l2(59),coll_y_l2(59),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(58),y_cood_l2(58),ball_x,ball_y,draw_l2(58),r_brick(58),g_brick(58),b_brick(58),coll_x_l2(58),coll_y_l2(58),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(57),y_cood_l2(57),ball_x,ball_y,draw_l2(57),r_brick(57),g_brick(57),b_brick(57),coll_x_l2(57),coll_y_l2(57),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(56),y_cood_l2(56),ball_x,ball_y,draw_l2(56),r_brick(56),g_brick(56),b_brick(56),coll_x_l2(56),coll_y_l2(56),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(55),y_cood_l2(55),ball_x,ball_y,draw_l2(55),r_brick(55),g_brick(55),b_brick(55),coll_x_l2(55),coll_y_l2(55),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(54),y_cood_l2(54),ball_x,ball_y,draw_l2(54),r_brick(54),g_brick(54),b_brick(54),coll_x_l2(54),coll_y_l2(54),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(53),y_cood_l2(53),ball_x,ball_y,draw_l2(53),r_brick(53),g_brick(53),b_brick(53),coll_x_l2(53),coll_y_l2(53),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(52),y_cood_l2(52),ball_x,ball_y,draw_l2(52),r_brick(52),g_brick(52),b_brick(52),coll_x_l2(52),coll_y_l2(52),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(51),y_cood_l2(51),ball_x,ball_y,draw_l2(51),r_brick(51),g_brick(51),b_brick(51),coll_x_l2(51),coll_y_l2(51),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(50),y_cood_l2(50),ball_x,ball_y,draw_l2(50),r_brick(50),g_brick(50),b_brick(50),coll_x_l2(50),coll_y_l2(50),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(49),y_cood_l2(49),ball_x,ball_y,draw_l2(49),r_brick(49),g_brick(49),b_brick(49),coll_x_l2(49),coll_y_l2(49),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(48),y_cood_l2(48),ball_x,ball_y,draw_l2(48),r_brick(48),g_brick(48),b_brick(48),coll_x_l2(48),coll_y_l2(48),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(47),y_cood_l2(47),ball_x,ball_y,draw_l2(47),r_brick(47),g_brick(47),b_brick(47),coll_x_l2(47),coll_y_l2(47),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(46),y_cood_l2(46),ball_x,ball_y,draw_l2(46),r_brick(46),g_brick(46),b_brick(46),coll_x_l2(46),coll_y_l2(46),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(45),y_cood_l2(45),ball_x,ball_y,draw_l2(45),r_brick(45),g_brick(45),b_brick(45),coll_x_l2(45),coll_y_l2(45),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l2(44),y_cood_l2(44),ball_x,ball_y,draw_l2(44),r_brick(44),g_brick(44),b_brick(44),coll_x_l2(44),coll_y_l2(44),ball_x_vel,ball_y_vel);	
							ball(hpos_scr,vpos_scr,ball_x,ball_y,ball_row,ball_col);	--get the ball image
						elsif(l3complete='0')then--display bricks of level 3
							brick(hpos_scr,vpos_scr,x_cood_l3(71),y_cood_l3(71),ball_x,ball_y,draw_l3(71),r_brick(71),g_brick(71),b_brick(71),coll_x_l3(71),coll_y_l3(71),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(70),y_cood_l3(70),ball_x,ball_y,draw_l3(70),r_brick(70),g_brick(70),b_brick(70),coll_x_l3(70),coll_y_l3(70),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(69),y_cood_l3(69),ball_x,ball_y,draw_l3(69),r_brick(69),g_brick(69),b_brick(69),coll_x_l3(69),coll_y_l3(69),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(68),y_cood_l3(68),ball_x,ball_y,draw_l3(68),r_brick(68),g_brick(68),b_brick(68),coll_x_l3(68),coll_y_l3(68),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(67),y_cood_l3(67),ball_x,ball_y,draw_l3(67),r_brick(67),g_brick(67),b_brick(67),coll_x_l3(67),coll_y_l3(67),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(66),y_cood_l3(66),ball_x,ball_y,draw_l3(66),r_brick(66),g_brick(66),b_brick(66),coll_x_l3(66),coll_y_l3(66),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(65),y_cood_l3(65),ball_x,ball_y,draw_l3(65),r_brick(65),g_brick(65),b_brick(65),coll_x_l3(65),coll_y_l3(65),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(64),y_cood_l3(64),ball_x,ball_y,draw_l3(64),r_brick(64),g_brick(64),b_brick(64),coll_x_l3(64),coll_y_l3(64),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(63),y_cood_l3(63),ball_x,ball_y,draw_l3(63),r_brick(63),g_brick(63),b_brick(63),coll_x_l3(63),coll_y_l3(63),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(62),y_cood_l3(62),ball_x,ball_y,draw_l3(62),r_brick(62),g_brick(62),b_brick(62),coll_x_l3(62),coll_y_l3(62),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(61),y_cood_l3(61),ball_x,ball_y,draw_l3(61),r_brick(61),g_brick(61),b_brick(61),coll_x_l3(61),coll_y_l3(61),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(60),y_cood_l3(60),ball_x,ball_y,draw_l3(60),r_brick(60),g_brick(60),b_brick(60),coll_x_l3(60),coll_y_l3(60),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(59),y_cood_l3(59),ball_x,ball_y,draw_l3(59),r_brick(59),g_brick(59),b_brick(59),coll_x_l3(59),coll_y_l3(59),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(58),y_cood_l3(58),ball_x,ball_y,draw_l3(58),r_brick(58),g_brick(58),b_brick(58),coll_x_l3(58),coll_y_l3(58),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(57),y_cood_l3(57),ball_x,ball_y,draw_l3(57),r_brick(57),g_brick(57),b_brick(57),coll_x_l3(57),coll_y_l3(57),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(56),y_cood_l3(56),ball_x,ball_y,draw_l3(56),r_brick(56),g_brick(56),b_brick(56),coll_x_l3(56),coll_y_l3(56),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(55),y_cood_l3(55),ball_x,ball_y,draw_l3(55),r_brick(55),g_brick(55),b_brick(55),coll_x_l3(55),coll_y_l3(55),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(54),y_cood_l3(54),ball_x,ball_y,draw_l3(54),r_brick(54),g_brick(54),b_brick(54),coll_x_l3(54),coll_y_l3(54),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(53),y_cood_l3(53),ball_x,ball_y,draw_l3(53),r_brick(53),g_brick(53),b_brick(53),coll_x_l3(53),coll_y_l3(53),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(52),y_cood_l3(52),ball_x,ball_y,draw_l3(52),r_brick(52),g_brick(52),b_brick(52),coll_x_l3(52),coll_y_l3(52),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(51),y_cood_l3(51),ball_x,ball_y,draw_l3(51),r_brick(51),g_brick(51),b_brick(51),coll_x_l3(51),coll_y_l3(51),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(50),y_cood_l3(50),ball_x,ball_y,draw_l3(50),r_brick(50),g_brick(50),b_brick(50),coll_x_l3(50),coll_y_l3(50),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(49),y_cood_l3(49),ball_x,ball_y,draw_l3(49),r_brick(49),g_brick(49),b_brick(49),coll_x_l3(49),coll_y_l3(49),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(48),y_cood_l3(48),ball_x,ball_y,draw_l3(48),r_brick(48),g_brick(48),b_brick(48),coll_x_l3(48),coll_y_l3(48),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(47),y_cood_l3(47),ball_x,ball_y,draw_l3(47),r_brick(47),g_brick(47),b_brick(47),coll_x_l3(47),coll_y_l3(47),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(46),y_cood_l3(46),ball_x,ball_y,draw_l3(46),r_brick(46),g_brick(46),b_brick(46),coll_x_l3(46),coll_y_l3(46),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(45),y_cood_l3(45),ball_x,ball_y,draw_l3(45),r_brick(45),g_brick(45),b_brick(45),coll_x_l3(45),coll_y_l3(45),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(44),y_cood_l3(44),ball_x,ball_y,draw_l3(44),r_brick(44),g_brick(44),b_brick(44),coll_x_l3(44),coll_y_l3(44),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(43),y_cood_l3(43),ball_x,ball_y,draw_l3(43),r_brick(43),g_brick(43),b_brick(43),coll_x_l3(43),coll_y_l3(43),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(42),y_cood_l3(42),ball_x,ball_y,draw_l3(42),r_brick(42),g_brick(42),b_brick(42),coll_x_l3(42),coll_y_l3(42),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(41),y_cood_l3(41),ball_x,ball_y,draw_l3(41),r_brick(41),g_brick(41),b_brick(41),coll_x_l3(41),coll_y_l3(41),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(40),y_cood_l3(40),ball_x,ball_y,draw_l3(40),r_brick(40),g_brick(40),b_brick(40),coll_x_l3(40),coll_y_l3(40),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(39),y_cood_l3(39),ball_x,ball_y,draw_l3(39),r_brick(39),g_brick(39),b_brick(39),coll_x_l3(39),coll_y_l3(39),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(38),y_cood_l3(38),ball_x,ball_y,draw_l3(38),r_brick(38),g_brick(38),b_brick(38),coll_x_l3(38),coll_y_l3(38),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(37),y_cood_l3(37),ball_x,ball_y,draw_l3(37),r_brick(37),g_brick(37),b_brick(37),coll_x_l3(37),coll_y_l3(37),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(36),y_cood_l3(36),ball_x,ball_y,draw_l3(36),r_brick(36),g_brick(36),b_brick(36),coll_x_l3(36),coll_y_l3(36),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(35),y_cood_l3(35),ball_x,ball_y,draw_l3(35),r_brick(35),g_brick(35),b_brick(35),coll_x_l3(35),coll_y_l3(35),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(34),y_cood_l3(34),ball_x,ball_y,draw_l3(34),r_brick(34),g_brick(34),b_brick(34),coll_x_l3(34),coll_y_l3(34),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(33),y_cood_l3(33),ball_x,ball_y,draw_l3(33),r_brick(33),g_brick(33),b_brick(33),coll_x_l3(33),coll_y_l3(33),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(32),y_cood_l3(32),ball_x,ball_y,draw_l3(32),r_brick(32),g_brick(32),b_brick(32),coll_x_l3(32),coll_y_l3(32),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(31),y_cood_l3(31),ball_x,ball_y,draw_l3(31),r_brick(31),g_brick(31),b_brick(31),coll_x_l3(31),coll_y_l3(31),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(30),y_cood_l3(30),ball_x,ball_y,draw_l3(30),r_brick(30),g_brick(30),b_brick(30),coll_x_l3(30),coll_y_l3(30),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(29),y_cood_l3(29),ball_x,ball_y,draw_l3(29),r_brick(29),g_brick(29),b_brick(29),coll_x_l3(29),coll_y_l3(29),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(28),y_cood_l3(28),ball_x,ball_y,draw_l3(28),r_brick(28),g_brick(28),b_brick(28),coll_x_l3(28),coll_y_l3(28),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(27),y_cood_l3(27),ball_x,ball_y,draw_l3(27),r_brick(27),g_brick(27),b_brick(27),coll_x_l3(27),coll_y_l3(27),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(26),y_cood_l3(26),ball_x,ball_y,draw_l3(26),r_brick(26),g_brick(26),b_brick(26),coll_x_l3(26),coll_y_l3(26),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(25),y_cood_l3(25),ball_x,ball_y,draw_l3(25),r_brick(25),g_brick(25),b_brick(25),coll_x_l3(25),coll_y_l3(25),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(24),y_cood_l3(24),ball_x,ball_y,draw_l3(24),r_brick(24),g_brick(24),b_brick(24),coll_x_l3(24),coll_y_l3(24),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(23),y_cood_l3(23),ball_x,ball_y,draw_l3(23),r_brick(23),g_brick(23),b_brick(23),coll_x_l3(23),coll_y_l3(23),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(22),y_cood_l3(22),ball_x,ball_y,draw_l3(22),r_brick(22),g_brick(22),b_brick(22),coll_x_l3(22),coll_y_l3(22),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(21),y_cood_l3(21),ball_x,ball_y,draw_l3(21),r_brick(21),g_brick(21),b_brick(21),coll_x_l3(21),coll_y_l3(21),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(20),y_cood_l3(20),ball_x,ball_y,draw_l3(20),r_brick(20),g_brick(20),b_brick(20),coll_x_l3(20),coll_y_l3(20),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(19),y_cood_l3(19),ball_x,ball_y,draw_l3(19),r_brick(19),g_brick(19),b_brick(19),coll_x_l3(19),coll_y_l3(19),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(18),y_cood_l3(18),ball_x,ball_y,draw_l3(18),r_brick(18),g_brick(18),b_brick(18),coll_x_l3(18),coll_y_l3(18),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(17),y_cood_l3(17),ball_x,ball_y,draw_l3(17),r_brick(17),g_brick(17),b_brick(17),coll_x_l3(17),coll_y_l3(17),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(16),y_cood_l3(16),ball_x,ball_y,draw_l3(16),r_brick(16),g_brick(16),b_brick(16),coll_x_l3(16),coll_y_l3(16),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(15),y_cood_l3(15),ball_x,ball_y,draw_l3(15),r_brick(15),g_brick(15),b_brick(15),coll_x_l3(15),coll_y_l3(15),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(14),y_cood_l3(14),ball_x,ball_y,draw_l3(14),r_brick(14),g_brick(14),b_brick(14),coll_x_l3(14),coll_y_l3(14),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(13),y_cood_l3(13),ball_x,ball_y,draw_l3(13),r_brick(13),g_brick(13),b_brick(13),coll_x_l3(13),coll_y_l3(13),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(12),y_cood_l3(12),ball_x,ball_y,draw_l3(12),r_brick(12),g_brick(12),b_brick(12),coll_x_l3(12),coll_y_l3(12),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(11),y_cood_l3(11),ball_x,ball_y,draw_l3(11),r_brick(11),g_brick(11),b_brick(11),coll_x_l3(11),coll_y_l3(11),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(10),y_cood_l3(10),ball_x,ball_y,draw_l3(10),r_brick(10),g_brick(10),b_brick(10),coll_x_l3(10),coll_y_l3(10),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(9),y_cood_l3(9),ball_x,ball_y,draw_l3(9),r_brick(9),g_brick(9),b_brick(9),coll_x_l3(9),coll_y_l3(9),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(8),y_cood_l3(8),ball_x,ball_y,draw_l3(8),r_brick(8),g_brick(8),b_brick(8),coll_x_l3(8),coll_y_l3(8),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(7),y_cood_l3(7),ball_x,ball_y,draw_l3(7),r_brick(7),g_brick(7),b_brick(7),coll_x_l3(7),coll_y_l3(7),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(6),y_cood_l3(6),ball_x,ball_y,draw_l3(6),r_brick(6),g_brick(6),b_brick(6),coll_x_l3(6),coll_y_l3(6),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(5),y_cood_l3(5),ball_x,ball_y,draw_l3(5),r_brick(5),g_brick(5),b_brick(5),coll_x_l3(5),coll_y_l3(5),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(4),y_cood_l3(4),ball_x,ball_y,draw_l3(4),r_brick(4),g_brick(4),b_brick(4),coll_x_l3(4),coll_y_l3(4),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(3),y_cood_l3(3),ball_x,ball_y,draw_l3(3),r_brick(3),g_brick(3),b_brick(3),coll_x_l3(3),coll_y_l3(3),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(2),y_cood_l3(2),ball_x,ball_y,draw_l3(2),r_brick(2),g_brick(2),b_brick(2),coll_x_l3(2),coll_y_l3(2),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(1),y_cood_l3(1),ball_x,ball_y,draw_l3(1),r_brick(1),g_brick(1),b_brick(1),coll_x_l3(1),coll_y_l3(1),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l3(0),y_cood_l3(0),ball_x,ball_y,draw_l3(0),r_brick(0),g_brick(0),b_brick(0),coll_x_l3(0),coll_y_l3(0),ball_x_vel,ball_y_vel);
						ball(hpos_scr,vpos_scr,ball_x,ball_y,ball_row,ball_col);	--get the ball image	
						elsif(l4complete='0')then--display bricks of level 4
							brick(hpos_scr,vpos_scr,x_cood_l4(71),y_cood_l4(71),ball_x,ball_y,draw_l4(71),r_brick(71),g_brick(71),b_brick(71),coll_x_l4(71),coll_y_l4(71),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(70),y_cood_l4(70),ball_x,ball_y,draw_l4(70),r_brick(70),g_brick(70),b_brick(70),coll_x_l4(70),coll_y_l4(70),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(69),y_cood_l4(69),ball_x,ball_y,draw_l4(69),r_brick(69),g_brick(69),b_brick(69),coll_x_l4(69),coll_y_l4(69),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(68),y_cood_l4(68),ball_x,ball_y,draw_l4(68),r_brick(68),g_brick(68),b_brick(68),coll_x_l4(68),coll_y_l4(68),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(67),y_cood_l4(67),ball_x,ball_y,draw_l4(67),r_brick(67),g_brick(67),b_brick(67),coll_x_l4(67),coll_y_l4(67),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(66),y_cood_l4(66),ball_x,ball_y,draw_l4(66),r_brick(66),g_brick(66),b_brick(66),coll_x_l4(66),coll_y_l4(66),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(65),y_cood_l4(65),ball_x,ball_y,draw_l4(65),r_brick(65),g_brick(65),b_brick(65),coll_x_l4(65),coll_y_l4(65),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(64),y_cood_l4(64),ball_x,ball_y,draw_l4(64),r_brick(64),g_brick(64),b_brick(64),coll_x_l4(64),coll_y_l4(64),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(63),y_cood_l4(63),ball_x,ball_y,draw_l4(63),r_brick(63),g_brick(63),b_brick(63),coll_x_l4(63),coll_y_l4(63),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(62),y_cood_l4(62),ball_x,ball_y,draw_l4(62),r_brick(62),g_brick(62),b_brick(62),coll_x_l4(62),coll_y_l4(62),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(61),y_cood_l4(61),ball_x,ball_y,draw_l4(61),r_brick(61),g_brick(61),b_brick(61),coll_x_l4(61),coll_y_l4(61),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(60),y_cood_l4(60),ball_x,ball_y,draw_l4(60),r_brick(60),g_brick(60),b_brick(60),coll_x_l4(60),coll_y_l4(60),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(59),y_cood_l4(59),ball_x,ball_y,draw_l4(59),r_brick(59),g_brick(59),b_brick(59),coll_x_l4(59),coll_y_l4(59),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(58),y_cood_l4(58),ball_x,ball_y,draw_l4(58),r_brick(58),g_brick(58),b_brick(58),coll_x_l4(58),coll_y_l4(58),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(57),y_cood_l4(57),ball_x,ball_y,draw_l4(57),r_brick(57),g_brick(57),b_brick(57),coll_x_l4(57),coll_y_l4(57),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(56),y_cood_l4(56),ball_x,ball_y,draw_l4(56),r_brick(56),g_brick(56),b_brick(56),coll_x_l4(56),coll_y_l4(56),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(55),y_cood_l4(55),ball_x,ball_y,draw_l4(55),r_brick(55),g_brick(55),b_brick(55),coll_x_l4(55),coll_y_l4(55),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(54),y_cood_l4(54),ball_x,ball_y,draw_l4(54),r_brick(54),g_brick(54),b_brick(54),coll_x_l4(54),coll_y_l4(54),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(53),y_cood_l4(53),ball_x,ball_y,draw_l4(53),r_brick(53),g_brick(53),b_brick(53),coll_x_l4(53),coll_y_l4(53),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(52),y_cood_l4(52),ball_x,ball_y,draw_l4(52),r_brick(52),g_brick(52),b_brick(52),coll_x_l4(52),coll_y_l4(52),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(51),y_cood_l4(51),ball_x,ball_y,draw_l4(51),r_brick(51),g_brick(51),b_brick(51),coll_x_l4(51),coll_y_l4(51),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(50),y_cood_l4(50),ball_x,ball_y,draw_l4(50),r_brick(50),g_brick(50),b_brick(50),coll_x_l4(50),coll_y_l4(50),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(49),y_cood_l4(49),ball_x,ball_y,draw_l4(49),r_brick(49),g_brick(49),b_brick(49),coll_x_l4(49),coll_y_l4(49),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(48),y_cood_l4(48),ball_x,ball_y,draw_l4(48),r_brick(48),g_brick(48),b_brick(48),coll_x_l4(48),coll_y_l4(48),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(47),y_cood_l4(47),ball_x,ball_y,draw_l4(47),r_brick(47),g_brick(47),b_brick(47),coll_x_l4(47),coll_y_l4(47),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(46),y_cood_l4(46),ball_x,ball_y,draw_l4(46),r_brick(46),g_brick(46),b_brick(46),coll_x_l4(46),coll_y_l4(46),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(45),y_cood_l4(45),ball_x,ball_y,draw_l4(45),r_brick(45),g_brick(45),b_brick(45),coll_x_l4(45),coll_y_l4(45),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(44),y_cood_l4(44),ball_x,ball_y,draw_l4(44),r_brick(44),g_brick(44),b_brick(44),coll_x_l4(44),coll_y_l4(44),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(43),y_cood_l4(43),ball_x,ball_y,draw_l4(43),r_brick(43),g_brick(43),b_brick(43),coll_x_l4(43),coll_y_l4(43),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(42),y_cood_l4(42),ball_x,ball_y,draw_l4(42),r_brick(42),g_brick(42),b_brick(42),coll_x_l4(42),coll_y_l4(42),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(41),y_cood_l4(41),ball_x,ball_y,draw_l4(41),r_brick(41),g_brick(41),b_brick(41),coll_x_l4(41),coll_y_l4(41),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(40),y_cood_l4(40),ball_x,ball_y,draw_l4(40),r_brick(40),g_brick(40),b_brick(40),coll_x_l4(40),coll_y_l4(40),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(39),y_cood_l4(39),ball_x,ball_y,draw_l4(39),r_brick(39),g_brick(39),b_brick(39),coll_x_l4(39),coll_y_l4(39),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(38),y_cood_l4(38),ball_x,ball_y,draw_l4(38),r_brick(38),g_brick(38),b_brick(38),coll_x_l4(38),coll_y_l4(38),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(37),y_cood_l4(37),ball_x,ball_y,draw_l4(37),r_brick(37),g_brick(37),b_brick(37),coll_x_l4(37),coll_y_l4(37),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(36),y_cood_l4(36),ball_x,ball_y,draw_l4(36),r_brick(36),g_brick(36),b_brick(36),coll_x_l4(36),coll_y_l4(36),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(35),y_cood_l4(35),ball_x,ball_y,draw_l4(35),r_brick(35),g_brick(35),b_brick(35),coll_x_l4(35),coll_y_l4(35),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(34),y_cood_l4(34),ball_x,ball_y,draw_l4(34),r_brick(34),g_brick(34),b_brick(34),coll_x_l4(34),coll_y_l4(34),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(33),y_cood_l4(33),ball_x,ball_y,draw_l4(33),r_brick(33),g_brick(33),b_brick(33),coll_x_l4(33),coll_y_l4(33),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(32),y_cood_l4(32),ball_x,ball_y,draw_l4(32),r_brick(32),g_brick(32),b_brick(32),coll_x_l4(32),coll_y_l4(32),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(31),y_cood_l4(31),ball_x,ball_y,draw_l4(31),r_brick(31),g_brick(31),b_brick(31),coll_x_l4(31),coll_y_l4(31),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(30),y_cood_l4(30),ball_x,ball_y,draw_l4(30),r_brick(30),g_brick(30),b_brick(30),coll_x_l4(30),coll_y_l4(30),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(29),y_cood_l4(29),ball_x,ball_y,draw_l4(29),r_brick(29),g_brick(29),b_brick(29),coll_x_l4(29),coll_y_l4(29),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(28),y_cood_l4(28),ball_x,ball_y,draw_l4(28),r_brick(28),g_brick(28),b_brick(28),coll_x_l4(28),coll_y_l4(28),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(27),y_cood_l4(27),ball_x,ball_y,draw_l4(27),r_brick(27),g_brick(27),b_brick(27),coll_x_l4(27),coll_y_l4(27),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(26),y_cood_l4(26),ball_x,ball_y,draw_l4(26),r_brick(26),g_brick(26),b_brick(26),coll_x_l4(26),coll_y_l4(26),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(25),y_cood_l4(25),ball_x,ball_y,draw_l4(25),r_brick(25),g_brick(25),b_brick(25),coll_x_l4(25),coll_y_l4(25),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(24),y_cood_l4(24),ball_x,ball_y,draw_l4(24),r_brick(24),g_brick(24),b_brick(24),coll_x_l4(24),coll_y_l4(24),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(23),y_cood_l4(23),ball_x,ball_y,draw_l4(23),r_brick(23),g_brick(23),b_brick(23),coll_x_l4(23),coll_y_l4(23),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(22),y_cood_l4(22),ball_x,ball_y,draw_l4(22),r_brick(22),g_brick(22),b_brick(22),coll_x_l4(22),coll_y_l4(22),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(21),y_cood_l4(21),ball_x,ball_y,draw_l4(21),r_brick(21),g_brick(21),b_brick(21),coll_x_l4(21),coll_y_l4(21),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(20),y_cood_l4(20),ball_x,ball_y,draw_l4(20),r_brick(20),g_brick(20),b_brick(20),coll_x_l4(20),coll_y_l4(20),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(19),y_cood_l4(19),ball_x,ball_y,draw_l4(19),r_brick(19),g_brick(19),b_brick(19),coll_x_l4(19),coll_y_l4(19),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(18),y_cood_l4(18),ball_x,ball_y,draw_l4(18),r_brick(18),g_brick(18),b_brick(18),coll_x_l4(18),coll_y_l4(18),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(17),y_cood_l4(17),ball_x,ball_y,draw_l4(17),r_brick(17),g_brick(17),b_brick(17),coll_x_l4(17),coll_y_l4(17),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(16),y_cood_l4(16),ball_x,ball_y,draw_l4(16),r_brick(16),g_brick(16),b_brick(16),coll_x_l4(16),coll_y_l4(16),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(15),y_cood_l4(15),ball_x,ball_y,draw_l4(15),r_brick(15),g_brick(15),b_brick(15),coll_x_l4(15),coll_y_l4(15),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(14),y_cood_l4(14),ball_x,ball_y,draw_l4(14),r_brick(14),g_brick(14),b_brick(14),coll_x_l4(14),coll_y_l4(14),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(13),y_cood_l4(13),ball_x,ball_y,draw_l4(13),r_brick(13),g_brick(13),b_brick(13),coll_x_l4(13),coll_y_l4(13),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(12),y_cood_l4(12),ball_x,ball_y,draw_l4(12),r_brick(12),g_brick(12),b_brick(12),coll_x_l4(12),coll_y_l4(12),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(11),y_cood_l4(11),ball_x,ball_y,draw_l4(11),r_brick(11),g_brick(11),b_brick(11),coll_x_l4(11),coll_y_l4(11),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(10),y_cood_l4(10),ball_x,ball_y,draw_l4(10),r_brick(10),g_brick(10),b_brick(10),coll_x_l4(10),coll_y_l4(10),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(9),y_cood_l4(9),ball_x,ball_y,draw_l4(9),r_brick(9),g_brick(9),b_brick(9),coll_x_l4(9),coll_y_l4(9),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l4(8),y_cood_l4(8),ball_x,ball_y,draw_l4(8),r_brick(8),g_brick(8),b_brick(8),coll_x_l4(8),coll_y_l4(8),ball_x_vel,ball_y_vel);
						ball(hpos_scr,vpos_scr,ball_x,ball_y,ball_row,ball_col);	--get the ball image	
						elsif(l5complete='0')then--display bricks of level 5
							brick(hpos_scr,vpos_scr,x_cood_l5(71),y_cood_l5(71),ball_x,ball_y,draw_l5(71),r_brick(71),g_brick(71),b_brick(71),coll_x_l5(71),coll_y_l5(71),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(70),y_cood_l5(70),ball_x,ball_y,draw_l5(70),r_brick(70),g_brick(70),b_brick(70),coll_x_l5(70),coll_y_l5(70),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(69),y_cood_l5(69),ball_x,ball_y,draw_l5(69),r_brick(69),g_brick(69),b_brick(69),coll_x_l5(69),coll_y_l5(69),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(68),y_cood_l5(68),ball_x,ball_y,draw_l5(68),r_brick(68),g_brick(68),b_brick(68),coll_x_l5(68),coll_y_l5(68),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(67),y_cood_l5(67),ball_x,ball_y,draw_l5(67),r_brick(67),g_brick(67),b_brick(67),coll_x_l5(67),coll_y_l5(67),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(66),y_cood_l5(66),ball_x,ball_y,draw_l5(66),r_brick(66),g_brick(66),b_brick(66),coll_x_l5(66),coll_y_l5(66),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(65),y_cood_l5(65),ball_x,ball_y,draw_l5(65),r_brick(65),g_brick(65),b_brick(65),coll_x_l5(65),coll_y_l5(65),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(64),y_cood_l5(64),ball_x,ball_y,draw_l5(64),r_brick(64),g_brick(64),b_brick(64),coll_x_l5(64),coll_y_l5(64),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(63),y_cood_l5(63),ball_x,ball_y,draw_l5(63),r_brick(63),g_brick(63),b_brick(63),coll_x_l5(63),coll_y_l5(63),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(62),y_cood_l5(62),ball_x,ball_y,draw_l5(62),r_brick(62),g_brick(62),b_brick(62),coll_x_l5(62),coll_y_l5(62),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(61),y_cood_l5(61),ball_x,ball_y,draw_l5(61),r_brick(61),g_brick(61),b_brick(61),coll_x_l5(61),coll_y_l5(61),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(60),y_cood_l5(60),ball_x,ball_y,draw_l5(60),r_brick(60),g_brick(60),b_brick(60),coll_x_l5(60),coll_y_l5(60),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(59),y_cood_l5(59),ball_x,ball_y,draw_l5(59),r_brick(59),g_brick(59),b_brick(59),coll_x_l5(59),coll_y_l5(59),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(58),y_cood_l5(58),ball_x,ball_y,draw_l5(58),r_brick(58),g_brick(58),b_brick(58),coll_x_l5(58),coll_y_l5(58),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(57),y_cood_l5(57),ball_x,ball_y,draw_l5(57),r_brick(57),g_brick(57),b_brick(57),coll_x_l5(57),coll_y_l5(57),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(56),y_cood_l5(56),ball_x,ball_y,draw_l5(56),r_brick(56),g_brick(56),b_brick(56),coll_x_l5(56),coll_y_l5(56),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(55),y_cood_l5(55),ball_x,ball_y,draw_l5(55),r_brick(55),g_brick(55),b_brick(55),coll_x_l5(55),coll_y_l5(55),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(54),y_cood_l5(54),ball_x,ball_y,draw_l5(54),r_brick(54),g_brick(54),b_brick(54),coll_x_l5(54),coll_y_l5(54),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(53),y_cood_l5(53),ball_x,ball_y,draw_l5(53),r_brick(53),g_brick(53),b_brick(53),coll_x_l5(53),coll_y_l5(53),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(52),y_cood_l5(52),ball_x,ball_y,draw_l5(52),r_brick(52),g_brick(52),b_brick(52),coll_x_l5(52),coll_y_l5(52),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(51),y_cood_l5(51),ball_x,ball_y,draw_l5(51),r_brick(51),g_brick(51),b_brick(51),coll_x_l5(51),coll_y_l5(51),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(50),y_cood_l5(50),ball_x,ball_y,draw_l5(50),r_brick(50),g_brick(50),b_brick(50),coll_x_l5(50),coll_y_l5(50),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(49),y_cood_l5(49),ball_x,ball_y,draw_l5(49),r_brick(49),g_brick(49),b_brick(49),coll_x_l5(49),coll_y_l5(49),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(48),y_cood_l5(48),ball_x,ball_y,draw_l5(48),r_brick(48),g_brick(48),b_brick(48),coll_x_l5(48),coll_y_l5(48),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(47),y_cood_l5(47),ball_x,ball_y,draw_l5(47),r_brick(47),g_brick(47),b_brick(47),coll_x_l5(47),coll_y_l5(47),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(46),y_cood_l5(46),ball_x,ball_y,draw_l5(46),r_brick(46),g_brick(46),b_brick(46),coll_x_l5(46),coll_y_l5(46),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(45),y_cood_l5(45),ball_x,ball_y,draw_l5(45),r_brick(45),g_brick(45),b_brick(45),coll_x_l5(45),coll_y_l5(45),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(44),y_cood_l5(44),ball_x,ball_y,draw_l5(44),r_brick(44),g_brick(44),b_brick(44),coll_x_l5(44),coll_y_l5(44),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(43),y_cood_l5(43),ball_x,ball_y,draw_l5(43),r_brick(43),g_brick(43),b_brick(43),coll_x_l5(43),coll_y_l5(43),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(42),y_cood_l5(42),ball_x,ball_y,draw_l5(42),r_brick(42),g_brick(42),b_brick(42),coll_x_l5(42),coll_y_l5(42),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(41),y_cood_l5(41),ball_x,ball_y,draw_l5(41),r_brick(41),g_brick(41),b_brick(41),coll_x_l5(41),coll_y_l5(41),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(40),y_cood_l5(40),ball_x,ball_y,draw_l5(40),r_brick(40),g_brick(40),b_brick(40),coll_x_l5(40),coll_y_l5(40),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(39),y_cood_l5(39),ball_x,ball_y,draw_l5(39),r_brick(39),g_brick(39),b_brick(39),coll_x_l5(39),coll_y_l5(39),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(38),y_cood_l5(38),ball_x,ball_y,draw_l5(38),r_brick(38),g_brick(38),b_brick(38),coll_x_l5(38),coll_y_l5(38),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(37),y_cood_l5(37),ball_x,ball_y,draw_l5(37),r_brick(37),g_brick(37),b_brick(37),coll_x_l5(37),coll_y_l5(37),ball_x_vel,ball_y_vel);
							brick(hpos_scr,vpos_scr,x_cood_l5(36),y_cood_l5(36),ball_x,ball_y,draw_l5(36),r_brick(36),g_brick(36),b_brick(36),coll_x_l5(36),coll_y_l5(36),ball_x_vel,ball_y_vel);
							ball(hpos_scr,vpos_scr,ball_x,ball_y,ball_row,ball_col);	--get the ball image
						else--all levels are completed sucessfully
							winmes(hpos_scr,vpos_scr,winmes_x,winmes_y,winmes_row,winmes_col);--get gameover image	
							stopball<='1';--to stop the ball motion
						end if;
						bat(hpos_scr,vpos_scr,bat_x,bat_y,draw_bat,r_bat,g_bat,b_bat);--display bat
						lives(hpos_scr,vpos_scr,lives_x,lives_y,lives_row,lives_col);--get lives image
					else--game has not started yet
						welmes(hpos_scr,vpos_scr,welmes_x,welmes_y,welmes_row,welmes_col);--welcome message
					end if;
					
					if(ball_y>480 and isalive=0) then--if last life is used uo
						gameover(hpos_scr,vpos_scr,gameover_x,gameover_y,gameover_row,gameover_col);--get gameover image		
						stopball<='1';--to stop the ball motion
					else
						null;
					end if;
					
					if(pause='1' and stopball='0' and notstarted='0')then--if pause switch is on
						paused(hpos_scr,vpos_scr,paused_x,paused_y,paused_row,paused_col);--get paused image			
					else
						null;
					end if;
					
				if(hpos>152 and hpos<793 and vpos>37 and vpos<518) then				
					if(welmes_validity_bit='1') then
						r<=r_welmes;	--display welcome message
						g<=g_welmes;
						b<=b_welmes;					
					elsif(lives_validity_bit='1') then
						r<=r_lives;	--display lives
						g<=g_lives;
						b<=b_lives;
					elsif(ball_validity_bit='1') then
						r<=r_ball;	--display ball
						g<=g_ball;
						b<=b_ball;
					elsif(draw_bat='1') then
						r<=r_bat;		--display bat
						g<=g_bat;
						b<=b_bat;
					elsif(paused_validity_bit='1') then
						r<=r_paused;	--display pause message
						g<=g_paused;
						b<=b_paused;
					elsif(gameover_validity_bit='1') then
						r<=r_gameover;	--display gameover
						g<=g_gameover;
						b<=b_gameover;	
					elsif(winmes_validity_bit='1') then
						r<=r_winmes;	--display winning message
						g<=g_winmes;
						b<=b_winmes;
					elsif(draw_l1(71)='1' and is_destroyed_l1(71)='0') then--display bricks of level1
						r<=r_brick(71);
						g<=g_brick(71);
						b<=b_brick(71);
					elsif(draw_l1(70)='1' and is_destroyed_l1(70)='0') then
						r<=r_brick(70);
						g<=g_brick(70);
						b<=b_brick(70);
					elsif(draw_l1(69)='1' and is_destroyed_l1(69)='0') then
						r<=r_brick(69);
						g<=g_brick(69);
						b<=b_brick(69);
					elsif(draw_l1(68)='1' and is_destroyed_l1(68)='0') then
						r<=r_brick(68);
						g<=g_brick(68);
						b<=b_brick(68);
					elsif(draw_l1(67)='1' and is_destroyed_l1(67)='0') then
						r<=r_brick(67);
						g<=g_brick(67);
						b<=b_brick(67);
					elsif(draw_l1(66)='1' and is_destroyed_l1(66)='0') then
						r<=r_brick(66);
						g<=g_brick(66);
						b<=b_brick(66);
					elsif(draw_l1(65)='1' and is_destroyed_l1(65)='0') then
						r<=r_brick(65);
						g<=g_brick(65);
						b<=b_brick(65);
					elsif(draw_l1(64)='1' and is_destroyed_l1(64)='0') then
						r<=r_brick(64);
						g<=g_brick(64);
						b<=b_brick(64);
						
					elsif(draw_l1(63)='1' and is_destroyed_l1(63)='0') then
						r<=r_brick(63);
						g<=g_brick(63);
						b<=b_brick(63);
					elsif(draw_l1(62)='1' and is_destroyed_l1(62)='0') then
						r<=r_brick(62);
						g<=g_brick(62);
						b<=b_brick(62);
					elsif(draw_l1(61)='1' and is_destroyed_l1(61)='0') then
						r<=r_brick(61);
						g<=g_brick(61);
						b<=b_brick(61);
					elsif(draw_l1(60)='1' and is_destroyed_l1(60)='0') then
						r<=r_brick(60);
						g<=g_brick(60);
						b<=b_brick(60);
					elsif(draw_l1(59)='1' and is_destroyed_l1(59)='0') then
						r<=r_brick(59);
						g<=g_brick(59);
						b<=b_brick(59);
					elsif(draw_l1(58)='1' and is_destroyed_l1(58)='0') then
						r<=r_brick(58);
						g<=g_brick(58);
						b<=b_brick(58);
					elsif(draw_l1(57)='1' and is_destroyed_l1(57)='0') then
						r<=r_brick(57);
						g<=g_brick(57);
						b<=b_brick(57);
					elsif(draw_l1(56)='1' and is_destroyed_l1(56)='0') then
						r<=r_brick(56);
						g<=g_brick(56);
						b<=b_brick(56);
						
					elsif(draw_l1(55)='1' and is_destroyed_l1(55)='0') then
						r<=r_brick(55);
						g<=g_brick(55);
						b<=b_brick(55);
					elsif(draw_l1(54)='1' and is_destroyed_l1(54)='0') then
						r<=r_brick(54);
						g<=g_brick(54);
						b<=b_brick(54);
					elsif(draw_l1(53)='1' and is_destroyed_l1(53)='0') then
						r<=r_brick(53);
						g<=g_brick(53);
						b<=b_brick(53);
					elsif(draw_l1(52)='1' and is_destroyed_l1(52)='0') then
						r<=r_brick(52);
						g<=g_brick(52);
						b<=b_brick(52);
					elsif(draw_l1(51)='1' and is_destroyed_l1(51)='0') then
						r<=r_brick(51);
						g<=g_brick(51);
						b<=b_brick(51);
					elsif(draw_l1(50)='1' and is_destroyed_l1(50)='0') then
						r<=r_brick(50);
						g<=g_brick(50);
						b<=b_brick(50);
					elsif(draw_l1(49)='1' and is_destroyed_l1(49)='0') then
						r<=r_brick(49);
						g<=g_brick(49);
						b<=b_brick(49);
					elsif(draw_l1(48)='1' and is_destroyed_l1(48)='0') then
						r<=r_brick(48);
						g<=g_brick(48);
						b<=b_brick(48);
						
					elsif(draw_l1(47)='1' and is_destroyed_l1(47)='0') then
						r<=r_brick(47);
						g<=g_brick(47);
						b<=b_brick(47);
					elsif(draw_l1(46)='1' and is_destroyed_l1(46)='0') then
						r<=r_brick(46);
						g<=g_brick(46);
						b<=b_brick(46);
					elsif(draw_l1(45)='1' and is_destroyed_l1(45)='0') then
						r<=r_brick(45);
						g<=g_brick(45);
						b<=b_brick(45);
					elsif(draw_l1(44)='1' and is_destroyed_l1(44)='0') then
						r<=r_brick(44);
						g<=g_brick(44);
						b<=b_brick(44);
					elsif(draw_l1(43)='1' and is_destroyed_l1(43)='0') then
						r<=r_brick(43);
						g<=g_brick(43);
						b<=b_brick(43);
					elsif(draw_l1(42)='1' and is_destroyed_l1(42)='0') then
						r<=r_brick(42);
						g<=g_brick(42);
						b<=b_brick(42);
					elsif(draw_l1(41)='1' and is_destroyed_l1(41)='0') then
						r<=r_brick(41);
						g<=g_brick(41);
						b<=b_brick(41);
					elsif(draw_l1(40)='1' and is_destroyed_l1(40)='0') then
						r<=r_brick(40);
						g<=g_brick(40);
						b<=b_brick(40);
						
					elsif(draw_l1(39)='1' and is_destroyed_l1(39)='0') then
						r<=r_brick(39);
						g<=g_brick(39);
						b<=b_brick(39);
					elsif(draw_l1(38)='1' and is_destroyed_l1(38)='0') then
						r<=r_brick(38);
						g<=g_brick(38);
						b<=b_brick(38);
					elsif(draw_l1(37)='1' and is_destroyed_l1(37)='0') then
						r<=r_brick(37);
						g<=g_brick(37);
						b<=b_brick(37);
					elsif(draw_l1(36)='1' and is_destroyed_l1(36)='0') then
						r<=r_brick(36);
						g<=g_brick(36);
						b<=b_brick(36);
					elsif(draw_l1(35)='1' and is_destroyed_l1(35)='0') then
						r<=r_brick(35);
						g<=g_brick(35);
						b<=b_brick(35);
					elsif(draw_l1(34)='1' and is_destroyed_l1(34)='0') then
						r<=r_brick(34);
						g<=g_brick(34);
						b<=b_brick(34);
					elsif(draw_l1(33)='1' and is_destroyed_l1(33)='0') then
						r<=r_brick(33);
						g<=g_brick(33);
						b<=b_brick(33);
					elsif(draw_l1(32)='1' and is_destroyed_l1(32)='0') then
						r<=r_brick(32);
						g<=g_brick(32);
						b<=b_brick(32);
						
					elsif(draw_l1(31)='1' and is_destroyed_l1(31)='0') then
						r<=r_brick(31);
						g<=g_brick(31);
						b<=b_brick(31);
					elsif(draw_l1(30)='1' and is_destroyed_l1(30)='0') then
						r<=r_brick(30);
						g<=g_brick(30);
						b<=b_brick(30);
					elsif(draw_l1(29)='1' and is_destroyed_l1(29)='0') then
						r<=r_brick(29);
						g<=g_brick(29);
						b<=b_brick(29);
					elsif(draw_l1(28)='1' and is_destroyed_l1(28)='0') then
						r<=r_brick(28);
						g<=g_brick(28);
						b<=b_brick(28);
					elsif(draw_l1(27)='1' and is_destroyed_l1(27)='0') then
						r<=r_brick(27);
						g<=g_brick(27);
						b<=b_brick(27);
					elsif(draw_l1(26)='1' and is_destroyed_l1(26)='0') then
						r<=r_brick(26);
						g<=g_brick(26);
						b<=b_brick(26);
					elsif(draw_l1(25)='1' and is_destroyed_l1(25)='0') then
						r<=r_brick(25);
						g<=g_brick(25);
						b<=b_brick(25);
					elsif(draw_l1(24)='1' and is_destroyed_l1(24)='0') then
						r<=r_brick(24);
						g<=g_brick(24);
						b<=b_brick(24);
						
					elsif(draw_l1(23)='1' and is_destroyed_l1(23)='0') then
						r<=r_brick(23);
						g<=g_brick(23);
						b<=b_brick(23);
					elsif(draw_l1(22)='1' and is_destroyed_l1(22)='0') then
						r<=r_brick(22);
						g<=g_brick(22);
						b<=b_brick(22);
					elsif(draw_l1(21)='1' and is_destroyed_l1(21)='0') then
						r<=r_brick(21);
						g<=g_brick(21);
						b<=b_brick(21);
					elsif(draw_l1(20)='1' and is_destroyed_l1(20)='0') then
						r<=r_brick(20);
						g<=g_brick(20);
						b<=b_brick(20);
					elsif(draw_l1(19)='1' and is_destroyed_l1(19)='0') then
						r<=r_brick(19);
						g<=g_brick(19);
						b<=b_brick(19);
					elsif(draw_l1(18)='1' and is_destroyed_l1(18)='0') then
						r<=r_brick(18);
						g<=g_brick(18);
						b<=b_brick(18);
					elsif(draw_l1(17)='1' and is_destroyed_l1(17)='0') then
						r<=r_brick(17);
						g<=g_brick(17);
						b<=b_brick(17);
					elsif(draw_l1(16)='1' and is_destroyed_l1(16)='0') then
						r<=r_brick(16);
						g<=g_brick(16);
						b<=b_brick(16);
						
					elsif(draw_l1(15)='1' and is_destroyed_l1(15)='0') then
						r<=r_brick(15);
						g<=g_brick(15);
						b<=b_brick(15);
					elsif(draw_l1(14)='1' and is_destroyed_l1(14)='0') then
						r<=r_brick(14);
						g<=g_brick(14);
						b<=b_brick(14);
					elsif(draw_l1(13)='1' and is_destroyed_l1(13)='0') then
						r<=r_brick(13);
						g<=g_brick(13);
						b<=b_brick(13);
					elsif(draw_l1(12)='1' and is_destroyed_l1(12)='0') then
						r<=r_brick(12);
						g<=g_brick(12);
						b<=b_brick(12);
					elsif(draw_l1(11)='1' and is_destroyed_l1(11)='0') then
						r<=r_brick(11);
						g<=g_brick(11);
						b<=b_brick(11);
					elsif(draw_l1(10)='1' and is_destroyed_l1(10)='0') then
						r<=r_brick(10);
						g<=g_brick(10);
						b<=b_brick(10);
					elsif(draw_l1(9)='1' and is_destroyed_l1(9)='0') then
						r<=r_brick(9);
						g<=g_brick(9);
						b<=b_brick(9);
					elsif(draw_l1(8)='1' and is_destroyed_l1(8)='0') then
						r<=r_brick(8);
						g<=g_brick(8);
						b<=b_brick(8);
						
					elsif(draw_l1(7)='1' and is_destroyed_l1(7)='0') then
						r<=r_brick(7);
						g<=g_brick(7);
						b<=b_brick(7);
					elsif(draw_l1(6)='1' and is_destroyed_l1(6)='0') then
						r<=r_brick(6);
						g<=g_brick(6);
						b<=b_brick(6);
					elsif(draw_l1(5)='1' and is_destroyed_l1(5)='0') then
						r<=r_brick(5);
						g<=g_brick(5);
						b<=b_brick(5);
					elsif(draw_l1(4)='1' and is_destroyed_l1(4)='0') then
						r<=r_brick(4);
						g<=g_brick(4);
						b<=b_brick(4);
					elsif(draw_l1(3)='1' and is_destroyed_l1(3)='0') then
						r<=r_brick(3);
						g<=g_brick(3);
						b<=b_brick(3);
					elsif(draw_l1(2)='1' and is_destroyed_l1(2)='0') then
						r<=r_brick(2);
						g<=g_brick(2);
						b<=b_brick(2);
					elsif(draw_l1(1)='1' and is_destroyed_l1(1)='0') then
						r<=r_brick(1);
						g<=g_brick(1);
						b<=b_brick(1);
					elsif(draw_l1(0)='1' and is_destroyed_l1(0)='0') then
						r<=r_brick(0);
						g<=g_brick(0);
						b<=b_brick(0);
						
					elsif(draw_l2(71)='1' and is_destroyed_l2(71)='0') then--display bricks of level2
						r<=r_brick(71);
						g<=g_brick(71);
						b<=b_brick(71);
					elsif(draw_l2(70)='1' and is_destroyed_l2(70)='0') then
						r<=r_brick(70);
						g<=g_brick(70);
						b<=b_brick(70);
					elsif(draw_l2(69)='1' and is_destroyed_l2(69)='0') then
						r<=r_brick(69);
						g<=g_brick(69);
						b<=b_brick(69);
					elsif(draw_l2(68)='1' and is_destroyed_l2(68)='0') then
						r<=r_brick(68);
						g<=g_brick(68);
						b<=b_brick(68);
					elsif(draw_l2(67)='1' and is_destroyed_l2(67)='0') then
						r<=r_brick(67);
						g<=g_brick(67);
						b<=b_brick(67);
					elsif(draw_l2(66)='1' and is_destroyed_l2(66)='0') then
						r<=r_brick(66);
						g<=g_brick(66);
						b<=b_brick(66);
					elsif(draw_l2(65)='1' and is_destroyed_l2(65)='0') then
						r<=r_brick(65);
						g<=g_brick(65);
						b<=b_brick(65);
					elsif(draw_l2(64)='1' and is_destroyed_l2(64)='0') then
						r<=r_brick(64);
						g<=g_brick(64);
						b<=b_brick(64);
						
					elsif(draw_l2(63)='1' and is_destroyed_l2(63)='0') then
						r<=r_brick(63);
						g<=g_brick(63);
						b<=b_brick(63);
					elsif(draw_l2(62)='1' and is_destroyed_l2(62)='0') then
						r<=r_brick(62);
						g<=g_brick(62);
						b<=b_brick(62);
					elsif(draw_l2(61)='1' and is_destroyed_l2(61)='0') then
						r<=r_brick(61);
						g<=g_brick(61);
						b<=b_brick(61);
					elsif(draw_l2(60)='1' and is_destroyed_l2(60)='0') then
						r<=r_brick(60);
						g<=g_brick(60);
						b<=b_brick(60);
					elsif(draw_l2(59)='1' and is_destroyed_l2(59)='0') then
						r<=r_brick(59);
						g<=g_brick(59);
						b<=b_brick(59);
					elsif(draw_l2(58)='1' and is_destroyed_l2(58)='0') then
						r<=r_brick(58);
						g<=g_brick(58);
						b<=b_brick(58);
					elsif(draw_l2(57)='1' and is_destroyed_l2(57)='0') then
						r<=r_brick(57);
						g<=g_brick(57);
						b<=b_brick(57);
					elsif(draw_l2(56)='1' and is_destroyed_l2(56)='0') then
						r<=r_brick(56);
						g<=g_brick(56);
						b<=b_brick(56);
						
					elsif(draw_l2(55)='1' and is_destroyed_l2(55)='0') then
						r<=r_brick(55);
						g<=g_brick(55);
						b<=b_brick(55);
					elsif(draw_l2(54)='1' and is_destroyed_l2(54)='0') then
						r<=r_brick(54);
						g<=g_brick(54);
						b<=b_brick(54);
					elsif(draw_l2(53)='1' and is_destroyed_l2(53)='0') then
						r<=r_brick(53);
						g<=g_brick(53);
						b<=b_brick(53);
					elsif(draw_l2(52)='1' and is_destroyed_l2(52)='0') then
						r<=r_brick(52);
						g<=g_brick(52);
						b<=b_brick(52);
					elsif(draw_l2(51)='1' and is_destroyed_l2(51)='0') then
						r<=r_brick(51);
						g<=g_brick(51);
						b<=b_brick(51);
					elsif(draw_l2(50)='1' and is_destroyed_l2(50)='0') then
						r<=r_brick(50);
						g<=g_brick(50);
						b<=b_brick(50);
					elsif(draw_l2(49)='1' and is_destroyed_l2(49)='0') then
						r<=r_brick(49);
						g<=g_brick(49);
						b<=b_brick(49);
					elsif(draw_l2(48)='1' and is_destroyed_l2(48)='0') then
						r<=r_brick(48);
						g<=g_brick(48);
						b<=b_brick(48);
						
					elsif(draw_l2(47)='1' and is_destroyed_l2(47)='0') then
						r<=r_brick(47);
						g<=g_brick(47);
						b<=b_brick(47);
					elsif(draw_l2(46)='1' and is_destroyed_l2(46)='0') then
						r<=r_brick(46);
						g<=g_brick(46);
						b<=b_brick(46);
					elsif(draw_l2(45)='1' and is_destroyed_l2(45)='0') then
						r<=r_brick(45);
						g<=g_brick(45);
						b<=b_brick(45);
					elsif(draw_l2(44)='1' and is_destroyed_l2(44)='0') then
						r<=r_brick(44);
						g<=g_brick(44);
						b<=b_brick(44);
						
					elsif(draw_l3(71)='1' and is_destroyed_l3(71)='0') then--display bricks of level3
						r<=r_brick(71);
						g<=g_brick(71);
						b<=b_brick(71);
					elsif(draw_l3(70)='1' and is_destroyed_l3(70)='0') then
						r<=r_brick(70);
						g<=g_brick(70);
						b<=b_brick(70);
					elsif(draw_l3(69)='1' and is_destroyed_l3(69)='0') then
						r<=r_brick(69);
						g<=g_brick(69);
						b<=b_brick(69);
					elsif(draw_l3(68)='1' and is_destroyed_l3(68)='0') then
						r<=r_brick(68);
						g<=g_brick(68);
						b<=b_brick(68);
					elsif(draw_l3(67)='1' and is_destroyed_l3(67)='0') then
						r<=r_brick(67);
						g<=g_brick(67);
						b<=b_brick(67);
					elsif(draw_l3(66)='1' and is_destroyed_l3(66)='0') then
						r<=r_brick(66);
						g<=g_brick(66);
						b<=b_brick(66);
					elsif(draw_l3(65)='1' and is_destroyed_l3(65)='0') then
						r<=r_brick(65);
						g<=g_brick(65);
						b<=b_brick(65);
					elsif(draw_l3(64)='1' and is_destroyed_l3(64)='0') then
						r<=r_brick(64);
						g<=g_brick(64);
						b<=b_brick(64);
						
					elsif(draw_l3(63)='1' and is_destroyed_l3(63)='0') then
						r<=r_brick(63);
						g<=g_brick(63);
						b<=b_brick(63);
					elsif(draw_l3(62)='1' and is_destroyed_l3(62)='0') then
						r<=r_brick(62);
						g<=g_brick(62);
						b<=b_brick(62);
					elsif(draw_l3(61)='1' and is_destroyed_l3(61)='0') then
						r<=r_brick(61);
						g<=g_brick(61);
						b<=b_brick(61);
					elsif(draw_l3(60)='1' and is_destroyed_l3(60)='0') then
						r<=r_brick(60);
						g<=g_brick(60);
						b<=b_brick(60);
					elsif(draw_l3(59)='1' and is_destroyed_l3(59)='0') then
						r<=r_brick(59);
						g<=g_brick(59);
						b<=b_brick(59);
					elsif(draw_l3(58)='1' and is_destroyed_l3(58)='0') then
						r<=r_brick(58);
						g<=g_brick(58);
						b<=b_brick(58);
					elsif(draw_l3(57)='1' and is_destroyed_l3(57)='0') then
						r<=r_brick(57);
						g<=g_brick(57);
						b<=b_brick(57);
					elsif(draw_l3(56)='1' and is_destroyed_l3(56)='0') then
						r<=r_brick(56);
						g<=g_brick(56);
						b<=b_brick(56);
						
					elsif(draw_l3(55)='1' and is_destroyed_l3(55)='0') then
						r<=r_brick(55);
						g<=g_brick(55);
						b<=b_brick(55);
					elsif(draw_l3(54)='1' and is_destroyed_l3(54)='0') then
						r<=r_brick(54);
						g<=g_brick(54);
						b<=b_brick(54);
					elsif(draw_l3(53)='1' and is_destroyed_l3(53)='0') then
						r<=r_brick(53);
						g<=g_brick(53);
						b<=b_brick(53);
					elsif(draw_l3(52)='1' and is_destroyed_l3(52)='0') then
						r<=r_brick(52);
						g<=g_brick(52);
						b<=b_brick(52);
					elsif(draw_l3(51)='1' and is_destroyed_l3(51)='0') then
						r<=r_brick(51);
						g<=g_brick(51);
						b<=b_brick(51);
					elsif(draw_l3(50)='1' and is_destroyed_l3(50)='0') then
						r<=r_brick(50);
						g<=g_brick(50);
						b<=b_brick(50);
					elsif(draw_l3(49)='1' and is_destroyed_l3(49)='0') then
						r<=r_brick(49);
						g<=g_brick(49);
						b<=b_brick(49);
					elsif(draw_l3(48)='1' and is_destroyed_l3(48)='0') then
						r<=r_brick(48);
						g<=g_brick(48);
						b<=b_brick(48);
						
					elsif(draw_l3(47)='1' and is_destroyed_l3(47)='0') then
						r<=r_brick(47);
						g<=g_brick(47);
						b<=b_brick(47);
					elsif(draw_l3(46)='1' and is_destroyed_l3(46)='0') then
						r<=r_brick(46);
						g<=g_brick(46);
						b<=b_brick(46);
					elsif(draw_l3(45)='1' and is_destroyed_l3(45)='0') then
						r<=r_brick(45);
						g<=g_brick(45);
						b<=b_brick(45);
					elsif(draw_l3(44)='1' and is_destroyed_l3(44)='0') then
						r<=r_brick(44);
						g<=g_brick(44);
						b<=b_brick(44);
					elsif(draw_l3(43)='1' and is_destroyed_l3(43)='0') then
						r<=r_brick(43);
						g<=g_brick(43);
						b<=b_brick(43);
					elsif(draw_l3(42)='1' and is_destroyed_l3(42)='0') then
						r<=r_brick(42);
						g<=g_brick(42);
						b<=b_brick(42);
					elsif(draw_l3(41)='1' and is_destroyed_l3(41)='0') then
						r<=r_brick(41);
						g<=g_brick(41);
						b<=b_brick(41);
					elsif(draw_l3(40)='1' and is_destroyed_l3(40)='0') then
						r<=r_brick(40);
						g<=g_brick(40);
						b<=b_brick(40);
						
					elsif(draw_l3(39)='1' and is_destroyed_l3(39)='0') then
						r<=r_brick(39);
						g<=g_brick(39);
						b<=b_brick(39);
					elsif(draw_l3(38)='1' and is_destroyed_l3(38)='0') then
						r<=r_brick(38);
						g<=g_brick(38);
						b<=b_brick(38);
					elsif(draw_l3(37)='1' and is_destroyed_l3(37)='0') then
						r<=r_brick(37);
						g<=g_brick(37);
						b<=b_brick(37);
					elsif(draw_l3(36)='1' and is_destroyed_l3(36)='0') then
						r<=r_brick(36);
						g<=g_brick(36);
						b<=b_brick(36);
					elsif(draw_l3(35)='1' and is_destroyed_l3(35)='0') then
						r<=r_brick(35);
						g<=g_brick(35);
						b<=b_brick(35);
					elsif(draw_l3(34)='1' and is_destroyed_l3(34)='0') then
						r<=r_brick(34);
						g<=g_brick(34);
						b<=b_brick(34);
					elsif(draw_l3(33)='1' and is_destroyed_l3(33)='0') then
						r<=r_brick(33);
						g<=g_brick(33);
						b<=b_brick(33);
					elsif(draw_l3(32)='1' and is_destroyed_l3(32)='0') then
						r<=r_brick(32);
						g<=g_brick(32);
						b<=b_brick(32);
						
					elsif(draw_l3(31)='1' and is_destroyed_l3(31)='0') then
						r<=r_brick(31);
						g<=g_brick(31);
						b<=b_brick(31);
					elsif(draw_l3(30)='1' and is_destroyed_l3(30)='0') then
						r<=r_brick(30);
						g<=g_brick(30);
						b<=b_brick(30);
					elsif(draw_l3(29)='1' and is_destroyed_l3(29)='0') then
						r<=r_brick(29);
						g<=g_brick(29);
						b<=b_brick(29);
					elsif(draw_l3(28)='1' and is_destroyed_l3(28)='0') then
						r<=r_brick(28);
						g<=g_brick(28);
						b<=b_brick(28);
					elsif(draw_l3(27)='1' and is_destroyed_l3(27)='0') then
						r<=r_brick(27);
						g<=g_brick(27);
						b<=b_brick(27);
					elsif(draw_l3(26)='1' and is_destroyed_l3(26)='0') then
						r<=r_brick(26);
						g<=g_brick(26);
						b<=b_brick(26);
					elsif(draw_l3(25)='1' and is_destroyed_l3(25)='0') then
						r<=r_brick(25);
						g<=g_brick(25);
						b<=b_brick(25);
					elsif(draw_l3(24)='1' and is_destroyed_l3(24)='0') then
						r<=r_brick(24);
						g<=g_brick(24);
						b<=b_brick(24);
						
					elsif(draw_l3(23)='1' and is_destroyed_l3(23)='0') then
						r<=r_brick(23);
						g<=g_brick(23);
						b<=b_brick(23);
					elsif(draw_l3(22)='1' and is_destroyed_l3(22)='0') then
						r<=r_brick(22);
						g<=g_brick(22);
						b<=b_brick(22);
					elsif(draw_l3(21)='1' and is_destroyed_l3(21)='0') then
						r<=r_brick(21);
						g<=g_brick(21);
						b<=b_brick(21);
					elsif(draw_l3(20)='1' and is_destroyed_l3(20)='0') then
						r<=r_brick(20);
						g<=g_brick(20);
						b<=b_brick(20);
					elsif(draw_l3(19)='1' and is_destroyed_l3(19)='0') then
						r<=r_brick(19);
						g<=g_brick(19);
						b<=b_brick(19);
					elsif(draw_l3(18)='1' and is_destroyed_l3(18)='0') then
						r<=r_brick(18);
						g<=g_brick(18);
						b<=b_brick(18);
					elsif(draw_l3(17)='1' and is_destroyed_l3(17)='0') then
						r<=r_brick(17);
						g<=g_brick(17);
						b<=b_brick(17);
					elsif(draw_l3(16)='1' and is_destroyed_l3(16)='0') then
						r<=r_brick(16);
						g<=g_brick(16);
						b<=b_brick(16);
						
					elsif(draw_l3(15)='1' and is_destroyed_l3(15)='0') then
						r<=r_brick(15);
						g<=g_brick(15);
						b<=b_brick(15);
					elsif(draw_l3(14)='1' and is_destroyed_l3(14)='0') then
						r<=r_brick(14);
						g<=g_brick(14);
						b<=b_brick(14);
					elsif(draw_l3(13)='1' and is_destroyed_l3(13)='0') then
						r<=r_brick(13);
						g<=g_brick(13);
						b<=b_brick(13);
					elsif(draw_l3(12)='1' and is_destroyed_l3(12)='0') then
						r<=r_brick(12);
						g<=g_brick(12);
						b<=b_brick(12);
					elsif(draw_l3(11)='1' and is_destroyed_l3(11)='0') then
						r<=r_brick(11);
						g<=g_brick(11);
						b<=b_brick(11);
					elsif(draw_l3(10)='1' and is_destroyed_l3(10)='0') then
						r<=r_brick(10);
						g<=g_brick(10);
						b<=b_brick(10);
					elsif(draw_l3(9)='1' and is_destroyed_l3(9)='0') then
						r<=r_brick(9);
						g<=g_brick(9);
						b<=b_brick(9);
					elsif(draw_l3(8)='1' and is_destroyed_l3(8)='0') then
						r<=r_brick(8);
						g<=g_brick(8);
						b<=b_brick(8);
						
					elsif(draw_l3(7)='1' and is_destroyed_l3(7)='0') then
						r<=r_brick(7);
						g<=g_brick(7);
						b<=b_brick(7);
					elsif(draw_l3(6)='1' and is_destroyed_l3(6)='0') then
						r<=r_brick(6);
						g<=g_brick(6);
						b<=b_brick(6);
					elsif(draw_l3(5)='1' and is_destroyed_l3(5)='0') then
						r<=r_brick(5);
						g<=g_brick(5);
						b<=b_brick(5);
					elsif(draw_l3(4)='1' and is_destroyed_l3(4)='0') then
						r<=r_brick(4);
						g<=g_brick(4);
						b<=b_brick(4);
					elsif(draw_l3(3)='1' and is_destroyed_l3(3)='0') then
						r<=r_brick(3);
						g<=g_brick(3);
						b<=b_brick(3);
					elsif(draw_l3(2)='1' and is_destroyed_l3(2)='0') then
						r<=r_brick(2);
						g<=g_brick(2);
						b<=b_brick(2);
					elsif(draw_l3(1)='1' and is_destroyed_l3(1)='0') then
						r<=r_brick(1);
						g<=g_brick(1);
						b<=b_brick(1);
					elsif(draw_l3(0)='1' and is_destroyed_l3(0)='0') then
						r<=r_brick(0);
						g<=g_brick(0);
						b<=b_brick(0);
															
					elsif(draw_l4(71)='1' and is_destroyed_l4(71)='0') then--display bricks of level4
						r<=r_brick(71);
						g<=g_brick(71);
						b<=b_brick(71);
					elsif(draw_l4(70)='1' and is_destroyed_l4(70)='0') then
						r<=r_brick(70);
						g<=g_brick(70);
						b<=b_brick(70);
					elsif(draw_l4(69)='1' and is_destroyed_l4(69)='0') then
						r<=r_brick(69);
						g<=g_brick(69);
						b<=b_brick(69);
					elsif(draw_l4(68)='1' and is_destroyed_l4(68)='0') then
						r<=r_brick(68);
						g<=g_brick(68);
						b<=b_brick(68);
					elsif(draw_l4(67)='1' and is_destroyed_l4(67)='0') then
						r<=r_brick(67);
						g<=g_brick(67);
						b<=b_brick(67);
					elsif(draw_l4(66)='1' and is_destroyed_l4(66)='0') then
						r<=r_brick(66);
						g<=g_brick(66);
						b<=b_brick(66);
					elsif(draw_l4(65)='1' and is_destroyed_l4(65)='0') then
						r<=r_brick(65);
						g<=g_brick(65);
						b<=b_brick(65);
					elsif(draw_l4(64)='1' and is_destroyed_l4(64)='0') then
						r<=r_brick(64);
						g<=g_brick(64);
						b<=b_brick(64);
						
					elsif(draw_l4(63)='1' and is_destroyed_l4(63)='0') then
						r<=r_brick(63);
						g<=g_brick(63);
						b<=b_brick(63);
					elsif(draw_l4(62)='1' and is_destroyed_l4(62)='0') then
						r<=r_brick(62);
						g<=g_brick(62);
						b<=b_brick(62);
					elsif(draw_l4(61)='1' and is_destroyed_l4(61)='0') then
						r<=r_brick(61);
						g<=g_brick(61);
						b<=b_brick(61);
					elsif(draw_l4(60)='1' and is_destroyed_l4(60)='0') then
						r<=r_brick(60);
						g<=g_brick(60);
						b<=b_brick(60);
					elsif(draw_l4(59)='1' and is_destroyed_l4(59)='0') then
						r<=r_brick(59);
						g<=g_brick(59);
						b<=b_brick(59);
					elsif(draw_l4(58)='1' and is_destroyed_l4(58)='0') then
						r<=r_brick(58);
						g<=g_brick(58);
						b<=b_brick(58);
					elsif(draw_l4(57)='1' and is_destroyed_l4(57)='0') then
						r<=r_brick(57);
						g<=g_brick(57);
						b<=b_brick(57);
					elsif(draw_l4(56)='1' and is_destroyed_l4(56)='0') then
						r<=r_brick(56);
						g<=g_brick(56);
						b<=b_brick(56);
						
					elsif(draw_l4(55)='1' and is_destroyed_l4(55)='0') then
						r<=r_brick(55);
						g<=g_brick(55);
						b<=b_brick(55);
					elsif(draw_l4(54)='1' and is_destroyed_l4(54)='0') then
						r<=r_brick(54);
						g<=g_brick(54);
						b<=b_brick(54);
					elsif(draw_l4(53)='1' and is_destroyed_l4(53)='0') then
						r<=r_brick(53);
						g<=g_brick(53);
						b<=b_brick(53);
					elsif(draw_l4(52)='1' and is_destroyed_l4(52)='0') then
						r<=r_brick(52);
						g<=g_brick(52);
						b<=b_brick(52);
					elsif(draw_l4(51)='1' and is_destroyed_l4(51)='0') then
						r<=r_brick(51);
						g<=g_brick(51);
						b<=b_brick(51);
					elsif(draw_l4(50)='1' and is_destroyed_l4(50)='0') then
						r<=r_brick(50);
						g<=g_brick(50);
						b<=b_brick(50);
					elsif(draw_l4(49)='1' and is_destroyed_l4(49)='0') then
						r<=r_brick(49);
						g<=g_brick(49);
						b<=b_brick(49);
					elsif(draw_l4(48)='1' and is_destroyed_l4(48)='0') then
						r<=r_brick(48);
						g<=g_brick(48);
						b<=b_brick(48);
						
					elsif(draw_l4(47)='1' and is_destroyed_l4(47)='0') then
						r<=r_brick(47);
						g<=g_brick(47);
						b<=b_brick(47);
					elsif(draw_l4(46)='1' and is_destroyed_l4(46)='0') then
						r<=r_brick(46);
						g<=g_brick(46);
						b<=b_brick(46);
					elsif(draw_l4(45)='1' and is_destroyed_l4(45)='0') then
						r<=r_brick(45);
						g<=g_brick(45);
						b<=b_brick(45);
					elsif(draw_l4(44)='1' and is_destroyed_l4(44)='0') then
						r<=r_brick(44);
						g<=g_brick(44);
						b<=b_brick(44);
					elsif(draw_l4(43)='1' and is_destroyed_l4(43)='0') then
						r<=r_brick(43);
						g<=g_brick(43);
						b<=b_brick(43);
					elsif(draw_l4(42)='1' and is_destroyed_l4(42)='0') then
						r<=r_brick(42);
						g<=g_brick(42);
						b<=b_brick(42);
					elsif(draw_l4(41)='1' and is_destroyed_l4(41)='0') then
						r<=r_brick(41);
						g<=g_brick(41);
						b<=b_brick(41);
					elsif(draw_l4(40)='1' and is_destroyed_l4(40)='0') then
						r<=r_brick(40);
						g<=g_brick(40);
						b<=b_brick(40);
						
					elsif(draw_l4(39)='1' and is_destroyed_l4(39)='0') then
						r<=r_brick(39);
						g<=g_brick(39);
						b<=b_brick(39);
					elsif(draw_l4(38)='1' and is_destroyed_l4(38)='0') then
						r<=r_brick(38);
						g<=g_brick(38);
						b<=b_brick(38);
					elsif(draw_l4(37)='1' and is_destroyed_l4(37)='0') then
						r<=r_brick(37);
						g<=g_brick(37);
						b<=b_brick(37);
					elsif(draw_l4(36)='1' and is_destroyed_l4(36)='0') then
						r<=r_brick(36);
						g<=g_brick(36);
						b<=b_brick(36);
					elsif(draw_l4(35)='1' and is_destroyed_l4(35)='0') then
						r<=r_brick(35);
						g<=g_brick(35);
						b<=b_brick(35);
					elsif(draw_l4(34)='1' and is_destroyed_l4(34)='0') then
						r<=r_brick(34);
						g<=g_brick(34);
						b<=b_brick(34);
					elsif(draw_l4(33)='1' and is_destroyed_l4(33)='0') then
						r<=r_brick(33);
						g<=g_brick(33);
						b<=b_brick(33);
					elsif(draw_l4(32)='1' and is_destroyed_l4(32)='0') then
						r<=r_brick(32);
						g<=g_brick(32);
						b<=b_brick(32);
						
					elsif(draw_l4(31)='1' and is_destroyed_l4(31)='0') then
						r<=r_brick(31);
						g<=g_brick(31);
						b<=b_brick(31);
					elsif(draw_l4(30)='1' and is_destroyed_l4(30)='0') then
						r<=r_brick(30);
						g<=g_brick(30);
						b<=b_brick(30);
					elsif(draw_l4(29)='1' and is_destroyed_l4(29)='0') then
						r<=r_brick(29);
						g<=g_brick(29);
						b<=b_brick(29);
					elsif(draw_l4(28)='1' and is_destroyed_l4(28)='0') then
						r<=r_brick(28);
						g<=g_brick(28);
						b<=b_brick(28);
					elsif(draw_l4(27)='1' and is_destroyed_l4(27)='0') then
						r<=r_brick(27);
						g<=g_brick(27);
						b<=b_brick(27);
					elsif(draw_l4(26)='1' and is_destroyed_l4(26)='0') then
						r<=r_brick(26);
						g<=g_brick(26);
						b<=b_brick(26);
					elsif(draw_l4(25)='1' and is_destroyed_l4(25)='0') then
						r<=r_brick(25);
						g<=g_brick(25);
						b<=b_brick(25);
					elsif(draw_l4(24)='1' and is_destroyed_l4(24)='0') then
						r<=r_brick(24);
						g<=g_brick(24);
						b<=b_brick(24);
						
					elsif(draw_l4(23)='1' and is_destroyed_l4(23)='0') then
						r<=r_brick(23);
						g<=g_brick(23);
						b<=b_brick(23);
					elsif(draw_l4(22)='1' and is_destroyed_l4(22)='0') then
						r<=r_brick(22);
						g<=g_brick(22);
						b<=b_brick(22);
					elsif(draw_l4(21)='1' and is_destroyed_l4(21)='0') then
						r<=r_brick(21);
						g<=g_brick(21);
						b<=b_brick(21);
					elsif(draw_l4(20)='1' and is_destroyed_l4(20)='0') then
						r<=r_brick(20);
						g<=g_brick(20);
						b<=b_brick(20);
					elsif(draw_l4(19)='1' and is_destroyed_l4(19)='0') then
						r<=r_brick(19);
						g<=g_brick(19);
						b<=b_brick(19);
					elsif(draw_l4(18)='1' and is_destroyed_l4(18)='0') then
						r<=r_brick(18);
						g<=g_brick(18);
						b<=b_brick(18);
					elsif(draw_l4(17)='1' and is_destroyed_l4(17)='0') then
						r<=r_brick(17);
						g<=g_brick(17);
						b<=b_brick(17);
					elsif(draw_l4(16)='1' and is_destroyed_l4(16)='0') then
						r<=r_brick(16);
						g<=g_brick(16);
						b<=b_brick(16);
						
					elsif(draw_l4(15)='1' and is_destroyed_l4(15)='0') then
						r<=r_brick(15);
						g<=g_brick(15);
						b<=b_brick(15);
					elsif(draw_l4(14)='1' and is_destroyed_l4(14)='0') then
						r<=r_brick(14);
						g<=g_brick(14);
						b<=b_brick(14);
					elsif(draw_l4(13)='1' and is_destroyed_l4(13)='0') then
						r<=r_brick(13);
						g<=g_brick(13);
						b<=b_brick(13);
					elsif(draw_l4(12)='1' and is_destroyed_l4(12)='0') then
						r<=r_brick(12);
						g<=g_brick(12);
						b<=b_brick(12);
					elsif(draw_l4(11)='1' and is_destroyed_l4(11)='0') then
						r<=r_brick(11);
						g<=g_brick(11);
						b<=b_brick(11);
					elsif(draw_l4(10)='1' and is_destroyed_l4(10)='0') then
						r<=r_brick(10);
						g<=g_brick(10);
						b<=b_brick(10);
					elsif(draw_l4(9)='1' and is_destroyed_l4(9)='0') then
						r<=r_brick(9);
						g<=g_brick(9);
						b<=b_brick(9);
					elsif(draw_l4(8)='1' and is_destroyed_l4(8)='0') then
						r<=r_brick(8);
						g<=g_brick(8);
						b<=b_brick(8);
						
					elsif(draw_l5(71)='1' and is_destroyed_l5(71)='0') then--display bricks of level5
						r<=r_brick(71);
						g<=g_brick(71);
						b<=b_brick(71);
					elsif(draw_l5(70)='1' and is_destroyed_l5(70)='0') then
						r<=r_brick(70);
						g<=g_brick(70);
						b<=b_brick(70);
					elsif(draw_l5(69)='1' and is_destroyed_l5(69)='0') then
						r<=r_brick(69);
						g<=g_brick(69);
						b<=b_brick(69);
					elsif(draw_l5(68)='1' and is_destroyed_l5(68)='0') then
						r<=r_brick(68);
						g<=g_brick(68);
						b<=b_brick(68);
					elsif(draw_l5(67)='1' and is_destroyed_l5(67)='0') then
						r<=r_brick(67);
						g<=g_brick(67);
						b<=b_brick(67);
					elsif(draw_l5(66)='1' and is_destroyed_l5(66)='0') then
						r<=r_brick(66);
						g<=g_brick(66);
						b<=b_brick(66);
					elsif(draw_l5(65)='1' and is_destroyed_l5(65)='0') then
						r<=r_brick(65);
						g<=g_brick(65);
						b<=b_brick(65);
					elsif(draw_l5(64)='1' and is_destroyed_l5(64)='0') then
						r<=r_brick(64);
						g<=g_brick(64);
						b<=b_brick(64);
						
					elsif(draw_l5(63)='1' and is_destroyed_l5(63)='0') then
						r<=r_brick(63);
						g<=g_brick(63);
						b<=b_brick(63);
					elsif(draw_l5(62)='1' and is_destroyed_l5(62)='0') then
						r<=r_brick(62);
						g<=g_brick(62);
						b<=b_brick(62);
					elsif(draw_l5(61)='1' and is_destroyed_l5(61)='0') then
						r<=r_brick(61);
						g<=g_brick(61);
						b<=b_brick(61);
					elsif(draw_l5(60)='1' and is_destroyed_l5(60)='0') then
						r<=r_brick(60);
						g<=g_brick(60);
						b<=b_brick(60);
					elsif(draw_l5(59)='1' and is_destroyed_l5(59)='0') then
						r<=r_brick(59);
						g<=g_brick(59);
						b<=b_brick(59);
					elsif(draw_l5(58)='1' and is_destroyed_l5(58)='0') then
						r<=r_brick(58);
						g<=g_brick(58);
						b<=b_brick(58);
					elsif(draw_l5(57)='1' and is_destroyed_l5(57)='0') then
						r<=r_brick(57);
						g<=g_brick(57);
						b<=b_brick(57);
					elsif(draw_l5(56)='1' and is_destroyed_l5(56)='0') then
						r<=r_brick(56);
						g<=g_brick(56);
						b<=b_brick(56);
						
					elsif(draw_l5(55)='1' and is_destroyed_l5(55)='0') then
						r<=r_brick(55);
						g<=g_brick(55);
						b<=b_brick(55);
					elsif(draw_l5(54)='1' and is_destroyed_l5(54)='0') then
						r<=r_brick(54);
						g<=g_brick(54);
						b<=b_brick(54);
					elsif(draw_l5(53)='1' and is_destroyed_l5(53)='0') then
						r<=r_brick(53);
						g<=g_brick(53);
						b<=b_brick(53);
					elsif(draw_l5(52)='1' and is_destroyed_l5(52)='0') then
						r<=r_brick(52);
						g<=g_brick(52);
						b<=b_brick(52);
					elsif(draw_l5(51)='1' and is_destroyed_l5(51)='0') then
						r<=r_brick(51);
						g<=g_brick(51);
						b<=b_brick(51);
					elsif(draw_l5(50)='1' and is_destroyed_l5(50)='0') then
						r<=r_brick(50);
						g<=g_brick(50);
						b<=b_brick(50);
					elsif(draw_l5(49)='1' and is_destroyed_l5(49)='0') then
						r<=r_brick(49);
						g<=g_brick(49);
						b<=b_brick(49);
					elsif(draw_l5(48)='1' and is_destroyed_l5(48)='0') then
						r<=r_brick(48);
						g<=g_brick(48);
						b<=b_brick(48);
						
					elsif(draw_l5(47)='1' and is_destroyed_l5(47)='0') then
						r<=r_brick(47);
						g<=g_brick(47);
						b<=b_brick(47);
					elsif(draw_l5(46)='1' and is_destroyed_l5(46)='0') then
						r<=r_brick(46);
						g<=g_brick(46);
						b<=b_brick(46);
					elsif(draw_l5(45)='1' and is_destroyed_l5(45)='0') then
						r<=r_brick(45);
						g<=g_brick(45);
						b<=b_brick(45);
					elsif(draw_l5(44)='1' and is_destroyed_l5(44)='0') then
						r<=r_brick(44);
						g<=g_brick(44);
						b<=b_brick(44);
					elsif(draw_l5(43)='1' and is_destroyed_l5(43)='0') then
						r<=r_brick(43);
						g<=g_brick(43);
						b<=b_brick(43);
					elsif(draw_l5(42)='1' and is_destroyed_l5(42)='0') then
						r<=r_brick(42);
						g<=g_brick(42);
						b<=b_brick(42);
					elsif(draw_l5(41)='1' and is_destroyed_l5(41)='0') then
						r<=r_brick(41);
						g<=g_brick(41);
						b<=b_brick(41);
					elsif(draw_l5(40)='1' and is_destroyed_l5(40)='0') then
						r<=r_brick(40);
						g<=g_brick(40);
						b<=b_brick(40);
						
					elsif(draw_l5(39)='1' and is_destroyed_l5(39)='0') then
						r<=r_brick(39);
						g<=g_brick(39);
						b<=b_brick(39);
					elsif(draw_l5(38)='1' and is_destroyed_l5(38)='0') then
						r<=r_brick(38);
						g<=g_brick(38);
						b<=b_brick(38);
					elsif(draw_l5(37)='1' and is_destroyed_l5(37)='0') then
						r<=r_brick(37);
						g<=g_brick(37);
						b<=b_brick(37);
					elsif(draw_l5(36)='1' and is_destroyed_l5(36)='0') then
						r<=r_brick(36);
						g<=g_brick(36);
						b<=b_brick(36);

					else
						r<="0000";	--if nothing then black screen
						g<="0000";
						b<="0000";
					end if;
				else
					r<="0000";	--make rgb 0 for period of fp,bp and sync duration
					g<="0000";
					b<="0000";
				end if;
					
					if(hpos<800) then
						hpos<=hpos+1;	--increment the horizontal pixel
					else
						hpos<=1;			--if entire line covered then reset
						if(vpos<525) then
							vpos<=vpos+1;	--increment the vertical pixel
						else
							vpos<=1;		--if entire screen covered then reset
								
							--1 means right direction or downwards
							--0 means left direction or upwards
							
							if(ball_x=5) then
								ball_x_vel<='1';	--if reached left edge then change direction to right
							elsif(ball_x=623) then
								ball_x_vel<='0';	--if reached right end then change direction to left
							else
								null;
							end if;
							
							if(ball_y=2) then
								ball_y_vel<='1';	--if reached top then reverse direction
							elsif(ball_y=448 and (ball_x>=bat_x-14 and ball_x<=bat_x+51)) then	--if reached bat height then check if hit the bat and then reverse direction else don't change
								ball_y_vel<='0';		
							else
								null;
							end if;
							
							if(is_destroyed_l1(71)='0')then--detect collision for ball and bricks of level1
								if(coll_x_l1(71)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(71)<='1';
								end if;
								if(coll_y_l1(71)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(71)<='1';
								end if;
							end if;
							if(is_destroyed_l1(70)='0')then
								if(coll_x_l1(70)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(70)<='1';
								end if;
								if(coll_y_l1(70)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(70)<='1';
								end if;
							end if;
							if(is_destroyed_l1(69)='0')then
								if(coll_x_l1(69)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(69)<='1';
								end if;
								if(coll_y_l1(69)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(69)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(68)='0')then
								if(coll_x_l1(68)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(68)<='1';
								end if;
								if(coll_y_l1(68)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(68)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(67)='0')then
								if(coll_x_l1(67)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(67)<='1';
								end if;
								if(coll_y_l1(67)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(67)<='1';
								end if;
							end if;
							if(is_destroyed_l1(66)='0')then
								if(coll_x_l1(66)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(66)<='1';
								end if;
								if(coll_y_l1(66)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(66)<='1';
								end if;
							end if;
							if(is_destroyed_l1(65)='0')then
								if(coll_x_l1(65)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(65)<='1';
								end if;
								if(coll_y_l1(65)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(65)<='1';
								end if;
							end if;
							if(is_destroyed_l1(64)='0')then
								if(coll_x_l1(64)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(64)<='1';
								end if;
								if(coll_y_l1(64)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(64)<='1';
								end if;
							end if;
							
							if(is_destroyed_l1(63)='0')then
								if(coll_x_l1(63)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(63)<='1';
								end if;
								if(coll_y_l1(63)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(63)<='1';
								end if;
							end if;
							if(is_destroyed_l1(62)='0')then
								if(coll_x_l1(62)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(62)<='1';
								end if;
								if(coll_y_l1(62)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(62)<='1';
								end if;
							end if;
							if(is_destroyed_l1(61)='0')then
								if(coll_x_l1(61)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(61)<='1';
								end if;
								if(coll_y_l1(61)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(61)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(60)='0')then
								if(coll_x_l1(60)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(60)<='1';
								end if;
								if(coll_y_l1(60)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(60)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(59)='0')then
								if(coll_x_l1(59)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(59)<='1';
								end if;
								if(coll_y_l1(59)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(59)<='1';
								end if;
							end if;
							if(is_destroyed_l1(58)='0')then
								if(coll_x_l1(58)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(58)<='1';
								end if;
								if(coll_y_l1(58)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(58)<='1';
								end if;
							end if;
							if(is_destroyed_l1(57)='0')then
								if(coll_x_l1(57)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(57)<='1';
								end if;
								if(coll_y_l1(57)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(57)<='1';
								end if;
							end if;
							if(is_destroyed_l1(56)='0')then
								if(coll_x_l1(56)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(56)<='1';
								end if;
								if(coll_y_l1(56)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(56)<='1';
								end if;
							end if;
							
							if(is_destroyed_l1(55)='0')then
								if(coll_x_l1(55)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(55)<='1';
								end if;
								if(coll_y_l1(55)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(55)<='1';
								end if;
							end if;
							if(is_destroyed_l1(54)='0')then
								if(coll_x_l1(54)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(54)<='1';
								end if;
								if(coll_y_l1(54)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(54)<='1';
								end if;
							end if;
							if(is_destroyed_l1(53)='0')then
								if(coll_x_l1(53)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(53)<='1';
								end if;
								if(coll_y_l1(53)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(53)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(52)='0')then
								if(coll_x_l1(52)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(52)<='1';
								end if;
								if(coll_y_l1(52)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(52)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(51)='0')then
								if(coll_x_l1(51)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(51)<='1';
								end if;
								if(coll_y_l1(51)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(51)<='1';
								end if;
							end if;
							if(is_destroyed_l1(50)='0')then
								if(coll_x_l1(50)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(50)<='1';
								end if;
								if(coll_y_l1(50)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(50)<='1';
								end if;
							end if;
							if(is_destroyed_l1(49)='0')then
								if(coll_x_l1(49)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(49)<='1';
								end if;
								if(coll_y_l1(49)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(49)<='1';
								end if;
							end if;
							if(is_destroyed_l1(48)='0')then
								if(coll_x_l1(48)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(48)<='1';
								end if;
								if(coll_y_l1(48)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(48)<='1';
								end if;
							end if;
							
							if(is_destroyed_l1(47)='0')then
								if(coll_x_l1(47)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(47)<='1';
								end if;
								if(coll_y_l1(47)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(47)<='1';
								end if;
							end if;
							if(is_destroyed_l1(46)='0')then
								if(coll_x_l1(46)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(46)<='1';
								end if;
								if(coll_y_l1(46)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(46)<='1';
								end if;
							end if;
							if(is_destroyed_l1(45)='0')then
								if(coll_x_l1(45)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(45)<='1';
								end if;
								if(coll_y_l1(45)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(45)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(44)='0')then
								if(coll_x_l1(44)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(44)<='1';
								end if;
								if(coll_y_l1(44)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(44)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(43)='0')then
								if(coll_x_l1(43)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(43)<='1';
								end if;
								if(coll_y_l1(43)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(43)<='1';
								end if;
							end if;
							if(is_destroyed_l1(42)='0')then
								if(coll_x_l1(42)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(42)<='1';
								end if;
								if(coll_y_l1(42)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(42)<='1';
								end if;
							end if;
							if(is_destroyed_l1(41)='0')then
								if(coll_x_l1(41)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(41)<='1';
								end if;
								if(coll_y_l1(41)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(41)<='1';
								end if;
							end if;
							if(is_destroyed_l1(40)='0')then
								if(coll_x_l1(40)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(40)<='1';
								end if;
								if(coll_y_l1(40)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(40)<='1';
								end if;
							end if;
							
							if(is_destroyed_l1(39)='0')then
								if(coll_x_l1(39)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(39)<='1';
								end if;
								if(coll_y_l1(39)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(39)<='1';
								end if;
							end if;
							if(is_destroyed_l1(38)='0')then
								if(coll_x_l1(38)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(38)<='1';
								end if;
								if(coll_y_l1(38)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(38)<='1';
								end if;
							end if;
							if(is_destroyed_l1(37)='0')then
								if(coll_x_l1(37)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(37)<='1';
								end if;
								if(coll_y_l1(37)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(37)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(36)='0')then
								if(coll_x_l1(36)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(36)<='1';
								end if;
								if(coll_y_l1(36)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(36)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(35)='0')then
								if(coll_x_l1(35)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(35)<='1';
								end if;
								if(coll_y_l1(35)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(35)<='1';
								end if;
							end if;
							if(is_destroyed_l1(34)='0')then
								if(coll_x_l1(34)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(34)<='1';
								end if;
								if(coll_y_l1(34)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(34)<='1';
								end if;
							end if;
							if(is_destroyed_l1(33)='0')then
								if(coll_x_l1(33)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(33)<='1';
								end if;
								if(coll_y_l1(33)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(33)<='1';
								end if;
							end if;
							if(is_destroyed_l1(32)='0')then
								if(coll_x_l1(32)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(32)<='1';
								end if;
								if(coll_y_l1(32)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(32)<='1';
								end if;
							end if;
							
							if(is_destroyed_l1(31)='0')then
								if(coll_x_l1(31)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(31)<='1';
								end if;
								if(coll_y_l1(31)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(31)<='1';
								end if;
							end if;
							if(is_destroyed_l1(30)='0')then
								if(coll_x_l1(30)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(30)<='1';
								end if;
								if(coll_y_l1(30)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(30)<='1';
								end if;
							end if;
							if(is_destroyed_l1(29)='0')then
								if(coll_x_l1(29)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(29)<='1';
								end if;
								if(coll_y_l1(29)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(29)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(28)='0')then
								if(coll_x_l1(28)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(28)<='1';
								end if;
								if(coll_y_l1(28)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(28)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(27)='0')then
								if(coll_x_l1(27)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(27)<='1';
								end if;
								if(coll_y_l1(27)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(27)<='1';
								end if;
							end if;
							if(is_destroyed_l1(26)='0')then
								if(coll_x_l1(26)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(26)<='1';
								end if;
								if(coll_y_l1(26)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(26)<='1';
								end if;
							end if;
							if(is_destroyed_l1(25)='0')then
								if(coll_x_l1(25)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(25)<='1';
								end if;
								if(coll_y_l1(25)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(25)<='1';
								end if;
							end if;
							if(is_destroyed_l1(24)='0')then
								if(coll_x_l1(24)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(24)<='1';
								end if;
								if(coll_y_l1(24)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(24)<='1';
								end if;
							end if;
							
							if(is_destroyed_l1(23)='0')then
								if(coll_x_l1(23)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(23)<='1';
								end if;
								if(coll_y_l1(23)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(23)<='1';
								end if;
							end if;
							if(is_destroyed_l1(22)='0')then
								if(coll_x_l1(22)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(22)<='1';
								end if;
								if(coll_y_l1(22)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(22)<='1';
								end if;
							end if;
							if(is_destroyed_l1(21)='0')then
								if(coll_x_l1(21)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(21)<='1';
								end if;
								if(coll_y_l1(21)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(21)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(20)='0')then
								if(coll_x_l1(20)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(20)<='1';
								end if;
								if(coll_y_l1(20)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(20)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(19)='0')then
								if(coll_x_l1(19)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(19)<='1';
								end if;
								if(coll_y_l1(19)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(19)<='1';
								end if;
							end if;
							if(is_destroyed_l1(18)='0')then
								if(coll_x_l1(18)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(18)<='1';
								end if;
								if(coll_y_l1(18)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(18)<='1';
								end if;
							end if;
							if(is_destroyed_l1(17)='0')then
								if(coll_x_l1(17)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(17)<='1';
								end if;
								if(coll_y_l1(17)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(17)<='1';
								end if;
							end if;
							if(is_destroyed_l1(16)='0')then
								if(coll_x_l1(16)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(16)<='1';
								end if;
								if(coll_y_l1(16)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(16)<='1';
								end if;
							end if;
							
							if(is_destroyed_l1(15)='0')then
								if(coll_x_l1(15)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(15)<='1';
								end if;
								if(coll_y_l1(15)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(15)<='1';
								end if;
							end if;
							if(is_destroyed_l1(14)='0')then
								if(coll_x_l1(14)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(14)<='1';
								end if;
								if(coll_y_l1(14)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(14)<='1';
								end if;
							end if;
							if(is_destroyed_l1(13)='0')then
								if(coll_x_l1(13)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(13)<='1';
								end if;
								if(coll_y_l1(13)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(13)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(12)='0')then
								if(coll_x_l1(12)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(12)<='1';
								end if;
								if(coll_y_l1(12)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(12)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(11)='0')then
								if(coll_x_l1(11)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(11)<='1';
								end if;
								if(coll_y_l1(11)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(11)<='1';
								end if;
							end if;
							if(is_destroyed_l1(10)='0')then
								if(coll_x_l1(10)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(10)<='1';
								end if;
								if(coll_y_l1(10)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(10)<='1';
								end if;
							end if;
							if(is_destroyed_l1(9)='0')then
								if(coll_x_l1(9)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(9)<='1';
								end if;
								if(coll_y_l1(9)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(9)<='1';
								end if;
							end if;
							if(is_destroyed_l1(8)='0')then
								if(coll_x_l1(8)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(8)<='1';
								end if;
								if(coll_y_l1(8)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(8)<='1';
								end if;
							end if;
							
							if(is_destroyed_l1(7)='0')then
								if(coll_x_l1(7)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(7)<='1';
								end if;
								if(coll_y_l1(7)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(7)<='1';
								end if;
							end if;
							if(is_destroyed_l1(6)='0')then
								if(coll_x_l1(6)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(6)<='1';
								end if;
								if(coll_y_l1(6)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(6)<='1';
								end if;
							end if;
							if(is_destroyed_l1(5)='0')then
								if(coll_x_l1(5)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(5)<='1';
								end if;
								if(coll_y_l1(5)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(5)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(4)='0')then
								if(coll_x_l1(4)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(4)<='1';
								end if;
								if(coll_y_l1(4)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(4)<='1';
								end if;
							end if;						
							if(is_destroyed_l1(3)='0')then
								if(coll_x_l1(3)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(3)<='1';
								end if;
								if(coll_y_l1(3)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(3)<='1';
								end if;
							end if;
							if(is_destroyed_l1(2)='0')then
								if(coll_x_l1(2)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(2)<='1';
								end if;
								if(coll_y_l1(2)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(2)<='1';
								end if;
							end if;
							if(is_destroyed_l1(1)='0')then
								if(coll_x_l1(1)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(1)<='1';
								end if;
								if(coll_y_l1(1)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(1)<='1';
								end if;
							end if;
							if(is_destroyed_l1(0)='0')then
								if(coll_x_l1(0)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l1(0)<='1';
								end if;
								if(coll_y_l1(0)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l1(0)<='1';
								end if;
							end if;
							
							if(is_destroyed_l2(71)='0')then--detect collision for ball and bricks of level2
								if(coll_x_l2(71)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(71)<='1';
								end if;
								if(coll_y_l2(71)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(71)<='1';
								end if;
							end if;
							if(is_destroyed_l2(70)='0')then
								if(coll_x_l2(70)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(70)<='1';
								end if;
								if(coll_y_l2(70)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(70)<='1';
								end if;
							end if;
							if(is_destroyed_l2(69)='0')then
								if(coll_x_l2(69)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(69)<='1';
								end if;
								if(coll_y_l2(69)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(69)<='1';
								end if;
							end if;						
							if(is_destroyed_l2(68)='0')then
								if(coll_x_l2(68)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(68)<='1';
								end if;
								if(coll_y_l2(68)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(68)<='1';
								end if;
							end if;						
							if(is_destroyed_l2(67)='0')then
								if(coll_x_l2(67)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(67)<='1';
								end if;
								if(coll_y_l2(67)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(67)<='1';
								end if;
							end if;
							if(is_destroyed_l2(66)='0')then
								if(coll_x_l2(66)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(66)<='1';
								end if;
								if(coll_y_l2(66)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(66)<='1';
								end if;
							end if;
							if(is_destroyed_l2(65)='0')then
								if(coll_x_l2(65)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(65)<='1';
								end if;
								if(coll_y_l2(65)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(65)<='1';
								end if;
							end if;
							if(is_destroyed_l2(64)='0')then
								if(coll_x_l2(64)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(64)<='1';
								end if;
								if(coll_y_l2(64)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(64)<='1';
								end if;
							end if;
							
							if(is_destroyed_l2(63)='0')then
								if(coll_x_l2(63)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(63)<='1';
								end if;
								if(coll_y_l2(63)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(63)<='1';
								end if;
							end if;
							if(is_destroyed_l2(62)='0')then
								if(coll_x_l2(62)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(62)<='1';
								end if;
								if(coll_y_l2(62)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(62)<='1';
								end if;
							end if;
							if(is_destroyed_l2(61)='0')then
								if(coll_x_l2(61)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(61)<='1';
								end if;
								if(coll_y_l2(61)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(61)<='1';
								end if;
							end if;						
							if(is_destroyed_l2(60)='0')then
								if(coll_x_l2(60)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(60)<='1';
								end if;
								if(coll_y_l2(60)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(60)<='1';
								end if;
							end if;						
							if(is_destroyed_l2(59)='0')then
								if(coll_x_l2(59)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(59)<='1';
								end if;
								if(coll_y_l2(59)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(59)<='1';
								end if;
							end if;
							if(is_destroyed_l2(58)='0')then
								if(coll_x_l2(58)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(58)<='1';
								end if;
								if(coll_y_l2(58)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(58)<='1';
								end if;
							end if;
							if(is_destroyed_l2(57)='0')then
								if(coll_x_l2(57)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(57)<='1';
								end if;
								if(coll_y_l2(57)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(57)<='1';
								end if;
							end if;
							if(is_destroyed_l2(56)='0')then
								if(coll_x_l2(56)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(56)<='1';
								end if;
								if(coll_y_l2(56)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(56)<='1';
								end if;
							end if;
							
							if(is_destroyed_l2(55)='0')then
								if(coll_x_l2(55)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(55)<='1';
								end if;
								if(coll_y_l2(55)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(55)<='1';
								end if;
							end if;
							if(is_destroyed_l2(54)='0')then
								if(coll_x_l2(54)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(54)<='1';
								end if;
								if(coll_y_l2(54)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(54)<='1';
								end if;
							end if;
							if(is_destroyed_l2(53)='0')then
								if(coll_x_l2(53)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(53)<='1';
								end if;
								if(coll_y_l2(53)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(53)<='1';
								end if;
							end if;						
							if(is_destroyed_l2(52)='0')then
								if(coll_x_l2(52)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(52)<='1';
								end if;
								if(coll_y_l2(52)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(52)<='1';
								end if;
							end if;						
							if(is_destroyed_l2(51)='0')then
								if(coll_x_l2(51)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(51)<='1';
								end if;
								if(coll_y_l2(51)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(51)<='1';
								end if;
							end if;
							if(is_destroyed_l2(50)='0')then
								if(coll_x_l2(50)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(50)<='1';
								end if;
								if(coll_y_l2(50)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(50)<='1';
								end if;
							end if;
							if(is_destroyed_l2(49)='0')then
								if(coll_x_l2(49)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(49)<='1';
								end if;
								if(coll_y_l2(49)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(49)<='1';
								end if;
							end if;
							if(is_destroyed_l2(48)='0')then
								if(coll_x_l2(48)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(48)<='1';
								end if;
								if(coll_y_l2(48)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(48)<='1';
								end if;
							end if;
							
							if(is_destroyed_l2(47)='0')then
								if(coll_x_l2(47)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(47)<='1';
								end if;
								if(coll_y_l2(47)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(47)<='1';
								end if;
							end if;
							if(is_destroyed_l2(46)='0')then
								if(coll_x_l2(46)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(46)<='1';
								end if;
								if(coll_y_l2(46)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(46)<='1';
								end if;
							end if;
							if(is_destroyed_l2(45)='0')then
								if(coll_x_l2(45)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(45)<='1';
								end if;
								if(coll_y_l2(45)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(45)<='1';
								end if;
							end if;						
							if(is_destroyed_l2(44)='0')then
								if(coll_x_l2(44)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l2(44)<='1';
								end if;
								if(coll_y_l2(44)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l2(44)<='1';
								end if;
							end if;
							
							if(is_destroyed_l3(71)='0')then--detect collision for ball and bricks of level3
								if(coll_x_l3(71)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(71)<='1';
								end if;
								if(coll_y_l3(71)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(71)<='1';
								end if;
							end if;
							if(is_destroyed_l3(70)='0')then
								if(coll_x_l3(70)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(70)<='1';
								end if;
								if(coll_y_l3(70)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(70)<='1';
								end if;
							end if;
							if(is_destroyed_l3(69)='0')then
								if(coll_x_l3(69)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(69)<='1';
								end if;
								if(coll_y_l3(69)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(69)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(68)='0')then
								if(coll_x_l3(68)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(68)<='1';
								end if;
								if(coll_y_l3(68)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(68)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(67)='0')then
								if(coll_x_l3(67)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(67)<='1';
								end if;
								if(coll_y_l3(67)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(67)<='1';
								end if;
							end if;
							if(is_destroyed_l3(66)='0')then
								if(coll_x_l3(66)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(66)<='1';
								end if;
								if(coll_y_l3(66)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(66)<='1';
								end if;
							end if;
							if(is_destroyed_l3(65)='0')then
								if(coll_x_l3(65)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(65)<='1';
								end if;
								if(coll_y_l3(65)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(65)<='1';
								end if;
							end if;
							if(is_destroyed_l3(64)='0')then
								if(coll_x_l3(64)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(64)<='1';
								end if;
								if(coll_y_l3(64)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(64)<='1';
								end if;
							end if;
							
							if(is_destroyed_l3(63)='0')then
								if(coll_x_l3(63)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(63)<='1';
								end if;
								if(coll_y_l3(63)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(63)<='1';
								end if;
							end if;
							if(is_destroyed_l3(62)='0')then
								if(coll_x_l3(62)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(62)<='1';
								end if;
								if(coll_y_l3(62)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(62)<='1';
								end if;
							end if;
							if(is_destroyed_l3(61)='0')then
								if(coll_x_l3(61)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(61)<='1';
								end if;
								if(coll_y_l3(61)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(61)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(60)='0')then
								if(coll_x_l3(60)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(60)<='1';
								end if;
								if(coll_y_l3(60)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(60)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(59)='0')then
								if(coll_x_l3(59)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(59)<='1';
								end if;
								if(coll_y_l3(59)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(59)<='1';
								end if;
							end if;
							if(is_destroyed_l3(58)='0')then
								if(coll_x_l3(58)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(58)<='1';
								end if;
								if(coll_y_l3(58)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(58)<='1';
								end if;
							end if;
							if(is_destroyed_l3(57)='0')then
								if(coll_x_l3(57)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(57)<='1';
								end if;
								if(coll_y_l3(57)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(57)<='1';
								end if;
							end if;
							if(is_destroyed_l3(56)='0')then
								if(coll_x_l3(56)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(56)<='1';
								end if;
								if(coll_y_l3(56)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(56)<='1';
								end if;
							end if;
							
							if(is_destroyed_l3(55)='0')then
								if(coll_x_l3(55)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(55)<='1';
								end if;
								if(coll_y_l3(55)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(55)<='1';
								end if;
							end if;
							if(is_destroyed_l3(54)='0')then
								if(coll_x_l3(54)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(54)<='1';
								end if;
								if(coll_y_l3(54)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(54)<='1';
								end if;
							end if;
							if(is_destroyed_l3(53)='0')then
								if(coll_x_l3(53)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(53)<='1';
								end if;
								if(coll_y_l3(53)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(53)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(52)='0')then
								if(coll_x_l3(52)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(52)<='1';
								end if;
								if(coll_y_l3(52)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(52)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(51)='0')then
								if(coll_x_l3(51)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(51)<='1';
								end if;
								if(coll_y_l3(51)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(51)<='1';
								end if;
							end if;
							if(is_destroyed_l3(50)='0')then
								if(coll_x_l3(50)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(50)<='1';
								end if;
								if(coll_y_l3(50)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(50)<='1';
								end if;
							end if;
							if(is_destroyed_l3(49)='0')then
								if(coll_x_l3(49)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(49)<='1';
								end if;
								if(coll_y_l3(49)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(49)<='1';
								end if;
							end if;
							if(is_destroyed_l3(48)='0')then
								if(coll_x_l3(48)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(48)<='1';
								end if;
								if(coll_y_l3(48)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(48)<='1';
								end if;
							end if;
							
							if(is_destroyed_l3(47)='0')then
								if(coll_x_l3(47)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(47)<='1';
								end if;
								if(coll_y_l3(47)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(47)<='1';
								end if;
							end if;
							if(is_destroyed_l3(46)='0')then
								if(coll_x_l3(46)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(46)<='1';
								end if;
								if(coll_y_l3(46)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(46)<='1';
								end if;
							end if;
							if(is_destroyed_l3(45)='0')then
								if(coll_x_l3(45)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(45)<='1';
								end if;
								if(coll_y_l3(45)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(45)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(44)='0')then
								if(coll_x_l3(44)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(44)<='1';
								end if;
								if(coll_y_l3(44)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(44)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(43)='0')then
								if(coll_x_l3(43)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(43)<='1';
								end if;
								if(coll_y_l3(43)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(43)<='1';
								end if;
							end if;
							if(is_destroyed_l3(42)='0')then
								if(coll_x_l3(42)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(42)<='1';
								end if;
								if(coll_y_l3(42)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(42)<='1';
								end if;
							end if;
							if(is_destroyed_l3(41)='0')then
								if(coll_x_l3(41)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(41)<='1';
								end if;
								if(coll_y_l3(41)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(41)<='1';
								end if;
							end if;
							if(is_destroyed_l3(40)='0')then
								if(coll_x_l3(40)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(40)<='1';
								end if;
								if(coll_y_l3(40)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(40)<='1';
								end if;
							end if;
							
							if(is_destroyed_l3(39)='0')then
								if(coll_x_l3(39)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(39)<='1';
								end if;
								if(coll_y_l3(39)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(39)<='1';
								end if;
							end if;
							if(is_destroyed_l3(38)='0')then
								if(coll_x_l3(38)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(38)<='1';
								end if;
								if(coll_y_l3(38)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(38)<='1';
								end if;
							end if;
							if(is_destroyed_l3(37)='0')then
								if(coll_x_l3(37)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(37)<='1';
								end if;
								if(coll_y_l3(37)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(37)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(36)='0')then
								if(coll_x_l3(36)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(36)<='1';
								end if;
								if(coll_y_l3(36)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(36)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(35)='0')then
								if(coll_x_l3(35)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(35)<='1';
								end if;
								if(coll_y_l3(35)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(35)<='1';
								end if;
							end if;
							if(is_destroyed_l3(34)='0')then
								if(coll_x_l3(34)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(34)<='1';
								end if;
								if(coll_y_l3(34)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(34)<='1';
								end if;
							end if;
							if(is_destroyed_l3(33)='0')then
								if(coll_x_l3(33)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(33)<='1';
								end if;
								if(coll_y_l3(33)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(33)<='1';
								end if;
							end if;
							if(is_destroyed_l3(32)='0')then
								if(coll_x_l3(32)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(32)<='1';
								end if;
								if(coll_y_l3(32)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(32)<='1';
								end if;
							end if;
							
							if(is_destroyed_l3(31)='0')then
								if(coll_x_l3(31)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(31)<='1';
								end if;
								if(coll_y_l3(31)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(31)<='1';
								end if;
							end if;
							if(is_destroyed_l3(30)='0')then
								if(coll_x_l3(30)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(30)<='1';
								end if;
								if(coll_y_l3(30)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(30)<='1';
								end if;
							end if;
							if(is_destroyed_l3(29)='0')then
								if(coll_x_l3(29)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(29)<='1';
								end if;
								if(coll_y_l3(29)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(29)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(28)='0')then
								if(coll_x_l3(28)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(28)<='1';
								end if;
								if(coll_y_l3(28)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(28)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(27)='0')then
								if(coll_x_l3(27)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(27)<='1';
								end if;
								if(coll_y_l3(27)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(27)<='1';
								end if;
							end if;
							if(is_destroyed_l3(26)='0')then
								if(coll_x_l3(26)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(26)<='1';
								end if;
								if(coll_y_l3(26)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(26)<='1';
								end if;
							end if;
							if(is_destroyed_l3(25)='0')then
								if(coll_x_l3(25)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(25)<='1';
								end if;
								if(coll_y_l3(25)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(25)<='1';
								end if;
							end if;
							if(is_destroyed_l3(24)='0')then
								if(coll_x_l3(24)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(24)<='1';
								end if;
								if(coll_y_l3(24)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(24)<='1';
								end if;
							end if;
							
							if(is_destroyed_l3(23)='0')then
								if(coll_x_l3(23)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(23)<='1';
								end if;
								if(coll_y_l3(23)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(23)<='1';
								end if;
							end if;
							if(is_destroyed_l3(22)='0')then
								if(coll_x_l3(22)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(22)<='1';
								end if;
								if(coll_y_l3(22)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(22)<='1';
								end if;
							end if;
							if(is_destroyed_l3(21)='0')then
								if(coll_x_l3(21)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(21)<='1';
								end if;
								if(coll_y_l3(21)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(21)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(20)='0')then
								if(coll_x_l3(20)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(20)<='1';
								end if;
								if(coll_y_l3(20)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(20)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(19)='0')then
								if(coll_x_l3(19)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(19)<='1';
								end if;
								if(coll_y_l3(19)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(19)<='1';
								end if;
							end if;
							if(is_destroyed_l3(18)='0')then
								if(coll_x_l3(18)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(18)<='1';
								end if;
								if(coll_y_l3(18)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(18)<='1';
								end if;
							end if;
							if(is_destroyed_l3(17)='0')then
								if(coll_x_l3(17)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(17)<='1';
								end if;
								if(coll_y_l3(17)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(17)<='1';
								end if;
							end if;
							if(is_destroyed_l3(16)='0')then
								if(coll_x_l3(16)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(16)<='1';
								end if;
								if(coll_y_l3(16)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(16)<='1';
								end if;
							end if;
							
							if(is_destroyed_l3(15)='0')then
								if(coll_x_l3(15)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(15)<='1';
								end if;
								if(coll_y_l3(15)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(15)<='1';
								end if;
							end if;
							if(is_destroyed_l3(14)='0')then
								if(coll_x_l3(14)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(14)<='1';
								end if;
								if(coll_y_l3(14)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(14)<='1';
								end if;
							end if;
							if(is_destroyed_l3(13)='0')then
								if(coll_x_l3(13)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(13)<='1';
								end if;
								if(coll_y_l3(13)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(13)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(12)='0')then
								if(coll_x_l3(12)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(12)<='1';
								end if;
								if(coll_y_l3(12)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(12)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(11)='0')then
								if(coll_x_l3(11)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(11)<='1';
								end if;
								if(coll_y_l3(11)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(11)<='1';
								end if;
							end if;
							if(is_destroyed_l3(10)='0')then
								if(coll_x_l3(10)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(10)<='1';
								end if;
								if(coll_y_l3(10)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(10)<='1';
								end if;
							end if;
							if(is_destroyed_l3(9)='0')then
								if(coll_x_l3(9)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(9)<='1';
								end if;
								if(coll_y_l3(9)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(9)<='1';
								end if;
							end if;
							if(is_destroyed_l3(8)='0')then
								if(coll_x_l3(8)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(8)<='1';
								end if;
								if(coll_y_l3(8)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(8)<='1';
								end if;
							end if;
							
							if(is_destroyed_l3(7)='0')then
								if(coll_x_l3(7)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(7)<='1';
								end if;
								if(coll_y_l3(7)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(7)<='1';
								end if;
							end if;
							if(is_destroyed_l3(6)='0')then
								if(coll_x_l3(6)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(6)<='1';
								end if;
								if(coll_y_l3(6)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(6)<='1';
								end if;
							end if;
							if(is_destroyed_l3(5)='0')then
								if(coll_x_l3(5)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(5)<='1';
								end if;
								if(coll_y_l3(5)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(5)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(4)='0')then
								if(coll_x_l3(4)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(4)<='1';
								end if;
								if(coll_y_l3(4)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(4)<='1';
								end if;
							end if;						
							if(is_destroyed_l3(3)='0')then
								if(coll_x_l3(3)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(3)<='1';
								end if;
								if(coll_y_l3(3)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(3)<='1';
								end if;
							end if;
							if(is_destroyed_l3(2)='0')then
								if(coll_x_l3(2)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(2)<='1';
								end if;
								if(coll_y_l3(2)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(2)<='1';
								end if;
							end if;
							if(is_destroyed_l3(1)='0')then
								if(coll_x_l3(1)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(1)<='1';
								end if;
								if(coll_y_l3(1)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(1)<='1';
								end if;
							end if;
							if(is_destroyed_l3(0)='0')then
								if(coll_x_l3(0)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l3(0)<='1';
								end if;
								if(coll_y_l3(0)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l3(0)<='1';
								end if;
							end if;
			
							if(is_destroyed_l4(71)='0')then--detect collision for ball and bricks of level4
								if(coll_x_l4(71)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(71)<='1';
								end if;
								if(coll_y_l4(71)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(71)<='1';
								end if;
							end if;
							if(is_destroyed_l4(70)='0')then
								if(coll_x_l4(70)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(70)<='1';
								end if;
								if(coll_y_l4(70)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(70)<='1';
								end if;
							end if;
							if(is_destroyed_l4(69)='0')then
								if(coll_x_l4(69)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(69)<='1';
								end if;
								if(coll_y_l4(69)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(69)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(68)='0')then
								if(coll_x_l4(68)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(68)<='1';
								end if;
								if(coll_y_l4(68)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(68)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(67)='0')then
								if(coll_x_l4(67)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(67)<='1';
								end if;
								if(coll_y_l4(67)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(67)<='1';
								end if;
							end if;
							if(is_destroyed_l4(66)='0')then
								if(coll_x_l4(66)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(66)<='1';
								end if;
								if(coll_y_l4(66)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(66)<='1';
								end if;
							end if;
							if(is_destroyed_l4(65)='0')then
								if(coll_x_l4(65)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(65)<='1';
								end if;
								if(coll_y_l4(65)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(65)<='1';
								end if;
							end if;
							if(is_destroyed_l4(64)='0')then
								if(coll_x_l4(64)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(64)<='1';
								end if;
								if(coll_y_l4(64)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(64)<='1';
								end if;
							end if;
							
							if(is_destroyed_l4(63)='0')then
								if(coll_x_l4(63)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(63)<='1';
								end if;
								if(coll_y_l4(63)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(63)<='1';
								end if;
							end if;
							if(is_destroyed_l4(62)='0')then
								if(coll_x_l4(62)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(62)<='1';
								end if;
								if(coll_y_l4(62)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(62)<='1';
								end if;
							end if;
							if(is_destroyed_l4(61)='0')then
								if(coll_x_l4(61)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(61)<='1';
								end if;
								if(coll_y_l4(61)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(61)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(60)='0')then
								if(coll_x_l4(60)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(60)<='1';
								end if;
								if(coll_y_l4(60)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(60)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(59)='0')then
								if(coll_x_l4(59)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(59)<='1';
								end if;
								if(coll_y_l4(59)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(59)<='1';
								end if;
							end if;
							if(is_destroyed_l4(58)='0')then
								if(coll_x_l4(58)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(58)<='1';
								end if;
								if(coll_y_l4(58)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(58)<='1';
								end if;
							end if;
							if(is_destroyed_l4(57)='0')then
								if(coll_x_l4(57)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(57)<='1';
								end if;
								if(coll_y_l4(57)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(57)<='1';
								end if;
							end if;
							if(is_destroyed_l4(56)='0')then
								if(coll_x_l4(56)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(56)<='1';
								end if;
								if(coll_y_l4(56)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(56)<='1';
								end if;
							end if;
							
							if(is_destroyed_l4(55)='0')then
								if(coll_x_l4(55)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(55)<='1';
								end if;
								if(coll_y_l4(55)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(55)<='1';
								end if;
							end if;
							if(is_destroyed_l4(54)='0')then
								if(coll_x_l4(54)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(54)<='1';
								end if;
								if(coll_y_l4(54)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(54)<='1';
								end if;
							end if;
							if(is_destroyed_l4(53)='0')then
								if(coll_x_l4(53)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(53)<='1';
								end if;
								if(coll_y_l4(53)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(53)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(52)='0')then
								if(coll_x_l4(52)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(52)<='1';
								end if;
								if(coll_y_l4(52)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(52)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(51)='0')then
								if(coll_x_l4(51)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(51)<='1';
								end if;
								if(coll_y_l4(51)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(51)<='1';
								end if;
							end if;
							if(is_destroyed_l4(50)='0')then
								if(coll_x_l4(50)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(50)<='1';
								end if;
								if(coll_y_l4(50)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(50)<='1';
								end if;
							end if;
							if(is_destroyed_l4(49)='0')then
								if(coll_x_l4(49)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(49)<='1';
								end if;
								if(coll_y_l4(49)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(49)<='1';
								end if;
							end if;
							if(is_destroyed_l4(48)='0')then
								if(coll_x_l4(48)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(48)<='1';
								end if;
								if(coll_y_l4(48)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(48)<='1';
								end if;
							end if;
							
							if(is_destroyed_l4(47)='0')then
								if(coll_x_l4(47)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(47)<='1';
								end if;
								if(coll_y_l4(47)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(47)<='1';
								end if;
							end if;
							if(is_destroyed_l4(46)='0')then
								if(coll_x_l4(46)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(46)<='1';
								end if;
								if(coll_y_l4(46)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(46)<='1';
								end if;
							end if;
							if(is_destroyed_l4(45)='0')then
								if(coll_x_l4(45)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(45)<='1';
								end if;
								if(coll_y_l4(45)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(45)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(44)='0')then
								if(coll_x_l4(44)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(44)<='1';
								end if;
								if(coll_y_l4(44)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(44)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(43)='0')then
								if(coll_x_l4(43)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(43)<='1';
								end if;
								if(coll_y_l4(43)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(43)<='1';
								end if;
							end if;
							if(is_destroyed_l4(42)='0')then
								if(coll_x_l4(42)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(42)<='1';
								end if;
								if(coll_y_l4(42)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(42)<='1';
								end if;
							end if;
							if(is_destroyed_l4(41)='0')then
								if(coll_x_l4(41)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(41)<='1';
								end if;
								if(coll_y_l4(41)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(41)<='1';
								end if;
							end if;
							if(is_destroyed_l4(40)='0')then
								if(coll_x_l4(40)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(40)<='1';
								end if;
								if(coll_y_l4(40)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(40)<='1';
								end if;
							end if;
							
							if(is_destroyed_l4(39)='0')then
								if(coll_x_l4(39)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(39)<='1';
								end if;
								if(coll_y_l4(39)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(39)<='1';
								end if;
							end if;
							if(is_destroyed_l4(38)='0')then
								if(coll_x_l4(38)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(38)<='1';
								end if;
								if(coll_y_l4(38)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(38)<='1';
								end if;
							end if;
							if(is_destroyed_l4(37)='0')then
								if(coll_x_l4(37)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(37)<='1';
								end if;
								if(coll_y_l4(37)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(37)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(36)='0')then
								if(coll_x_l4(36)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(36)<='1';
								end if;
								if(coll_y_l4(36)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(36)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(35)='0')then
								if(coll_x_l4(35)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(35)<='1';
								end if;
								if(coll_y_l4(35)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(35)<='1';
								end if;
							end if;
							if(is_destroyed_l4(34)='0')then
								if(coll_x_l4(34)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(34)<='1';
								end if;
								if(coll_y_l4(34)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(34)<='1';
								end if;
							end if;
							if(is_destroyed_l4(33)='0')then
								if(coll_x_l4(33)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(33)<='1';
								end if;
								if(coll_y_l4(33)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(33)<='1';
								end if;
							end if;
							if(is_destroyed_l4(32)='0')then
								if(coll_x_l4(32)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(32)<='1';
								end if;
								if(coll_y_l4(32)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(32)<='1';
								end if;
							end if;
							
							if(is_destroyed_l4(31)='0')then
								if(coll_x_l4(31)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(31)<='1';
								end if;
								if(coll_y_l4(31)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(31)<='1';
								end if;
							end if;
							if(is_destroyed_l4(30)='0')then
								if(coll_x_l4(30)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(30)<='1';
								end if;
								if(coll_y_l4(30)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(30)<='1';
								end if;
							end if;
							if(is_destroyed_l4(29)='0')then
								if(coll_x_l4(29)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(29)<='1';
								end if;
								if(coll_y_l4(29)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(29)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(28)='0')then
								if(coll_x_l4(28)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(28)<='1';
								end if;
								if(coll_y_l4(28)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(28)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(27)='0')then
								if(coll_x_l4(27)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(27)<='1';
								end if;
								if(coll_y_l4(27)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(27)<='1';
								end if;
							end if;
							if(is_destroyed_l4(26)='0')then
								if(coll_x_l4(26)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(26)<='1';
								end if;
								if(coll_y_l4(26)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(26)<='1';
								end if;
							end if;
							if(is_destroyed_l4(25)='0')then
								if(coll_x_l4(25)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(25)<='1';
								end if;
								if(coll_y_l4(25)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(25)<='1';
								end if;
							end if;
							if(is_destroyed_l4(24)='0')then
								if(coll_x_l4(24)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(24)<='1';
								end if;
								if(coll_y_l4(24)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(24)<='1';
								end if;
							end if;
							
							if(is_destroyed_l4(23)='0')then
								if(coll_x_l4(23)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(23)<='1';
								end if;
								if(coll_y_l4(23)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(23)<='1';
								end if;
							end if;
							if(is_destroyed_l4(22)='0')then
								if(coll_x_l4(22)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(22)<='1';
								end if;
								if(coll_y_l4(22)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(22)<='1';
								end if;
							end if;
							if(is_destroyed_l4(21)='0')then
								if(coll_x_l4(21)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(21)<='1';
								end if;
								if(coll_y_l4(21)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(21)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(20)='0')then
								if(coll_x_l4(20)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(20)<='1';
								end if;
								if(coll_y_l4(20)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(20)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(19)='0')then
								if(coll_x_l4(19)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(19)<='1';
								end if;
								if(coll_y_l4(19)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(19)<='1';
								end if;
							end if;
							if(is_destroyed_l4(18)='0')then
								if(coll_x_l4(18)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(18)<='1';
								end if;
								if(coll_y_l4(18)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(18)<='1';
								end if;
							end if;
							if(is_destroyed_l4(17)='0')then
								if(coll_x_l4(17)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(17)<='1';
								end if;
								if(coll_y_l4(17)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(17)<='1';
								end if;
							end if;
							if(is_destroyed_l4(16)='0')then
								if(coll_x_l4(16)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(16)<='1';
								end if;
								if(coll_y_l4(16)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(16)<='1';
								end if;
							end if;
							
							if(is_destroyed_l4(15)='0')then
								if(coll_x_l4(15)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(15)<='1';
								end if;
								if(coll_y_l4(15)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(15)<='1';
								end if;
							end if;
							if(is_destroyed_l4(14)='0')then
								if(coll_x_l4(14)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(14)<='1';
								end if;
								if(coll_y_l4(14)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(14)<='1';
								end if;
							end if;
							if(is_destroyed_l4(13)='0')then
								if(coll_x_l4(13)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(13)<='1';
								end if;
								if(coll_y_l4(13)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(13)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(12)='0')then
								if(coll_x_l4(12)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(12)<='1';
								end if;
								if(coll_y_l4(12)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(12)<='1';
								end if;
							end if;						
							if(is_destroyed_l4(11)='0')then
								if(coll_x_l4(11)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(11)<='1';
								end if;
								if(coll_y_l4(11)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(11)<='1';
								end if;
							end if;
							if(is_destroyed_l4(10)='0')then
								if(coll_x_l4(10)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(10)<='1';
								end if;
								if(coll_y_l4(10)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(10)<='1';
								end if;
							end if;
							if(is_destroyed_l4(9)='0')then
								if(coll_x_l4(9)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(9)<='1';
								end if;
								if(coll_y_l4(9)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(9)<='1';
								end if;
							end if;
							if(is_destroyed_l4(8)='0')then
								if(coll_x_l4(8)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l4(8)<='1';
								end if;
								if(coll_y_l4(8)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l4(8)<='1';
								end if;
							end if;
							
							if(is_destroyed_l5(71)='0')then--detect collision for ball and bricks of level5
								if(coll_x_l5(71)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(71)<='1';
								end if;
								if(coll_y_l5(71)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(71)<='1';
								end if;
							end if;
							if(is_destroyed_l5(70)='0')then
								if(coll_x_l5(70)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(70)<='1';
								end if;
								if(coll_y_l5(70)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(70)<='1';
								end if;
							end if;
							if(is_destroyed_l5(69)='0')then
								if(coll_x_l5(69)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(69)<='1';
								end if;
								if(coll_y_l5(69)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(69)<='1';
								end if;
							end if;						
							if(is_destroyed_l5(68)='0')then
								if(coll_x_l5(68)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(68)<='1';
								end if;
								if(coll_y_l5(68)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(68)<='1';
								end if;
							end if;						
							if(is_destroyed_l5(67)='0')then
								if(coll_x_l5(67)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(67)<='1';
								end if;
								if(coll_y_l5(67)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(67)<='1';
								end if;
							end if;
							if(is_destroyed_l5(66)='0')then
								if(coll_x_l5(66)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(66)<='1';
								end if;
								if(coll_y_l5(66)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(66)<='1';
								end if;
							end if;
							if(is_destroyed_l5(65)='0')then
								if(coll_x_l5(65)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(65)<='1';
								end if;
								if(coll_y_l5(65)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(65)<='1';
								end if;
							end if;
							if(is_destroyed_l5(64)='0')then
								if(coll_x_l5(64)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(64)<='1';
								end if;
								if(coll_y_l5(64)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(64)<='1';
								end if;
							end if;
							
							if(is_destroyed_l5(63)='0')then
								if(coll_x_l5(63)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(63)<='1';
								end if;
								if(coll_y_l5(63)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(63)<='1';
								end if;
							end if;
							if(is_destroyed_l5(62)='0')then
								if(coll_x_l5(62)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(62)<='1';
								end if;
								if(coll_y_l5(62)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(62)<='1';
								end if;
							end if;
							if(is_destroyed_l5(61)='0')then
								if(coll_x_l5(61)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(61)<='1';
								end if;
								if(coll_y_l5(61)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(61)<='1';
								end if;
							end if;						
							if(is_destroyed_l5(60)='0')then
								if(coll_x_l5(60)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(60)<='1';
								end if;
								if(coll_y_l5(60)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(60)<='1';
								end if;
							end if;						
							if(is_destroyed_l5(59)='0')then
								if(coll_x_l5(59)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(59)<='1';
								end if;
								if(coll_y_l5(59)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(59)<='1';
								end if;
							end if;
							if(is_destroyed_l5(58)='0')then
								if(coll_x_l5(58)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(58)<='1';
								end if;
								if(coll_y_l5(58)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(58)<='1';
								end if;
							end if;
							if(is_destroyed_l5(57)='0')then
								if(coll_x_l5(57)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(57)<='1';
								end if;
								if(coll_y_l5(57)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(57)<='1';
								end if;
							end if;
							if(is_destroyed_l5(56)='0')then
								if(coll_x_l5(56)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(56)<='1';
								end if;
								if(coll_y_l5(56)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(56)<='1';
								end if;
							end if;
							
							if(is_destroyed_l5(55)='0')then
								if(coll_x_l5(55)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(55)<='1';
								end if;
								if(coll_y_l5(55)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(55)<='1';
								end if;
							end if;
							if(is_destroyed_l5(54)='0')then
								if(coll_x_l5(54)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(54)<='1';
								end if;
								if(coll_y_l5(54)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(54)<='1';
								end if;
							end if;
							if(is_destroyed_l5(53)='0')then
								if(coll_x_l5(53)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(53)<='1';
								end if;
								if(coll_y_l5(53)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(53)<='1';
								end if;
							end if;						
							if(is_destroyed_l5(52)='0')then
								if(coll_x_l5(52)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(52)<='1';
								end if;
								if(coll_y_l5(52)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(52)<='1';
								end if;
							end if;						
							if(is_destroyed_l5(51)='0')then
								if(coll_x_l5(51)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(51)<='1';
								end if;
								if(coll_y_l5(51)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(51)<='1';
								end if;
							end if;
							if(is_destroyed_l5(50)='0')then
								if(coll_x_l5(50)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(50)<='1';
								end if;
								if(coll_y_l5(50)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(50)<='1';
								end if;
							end if;
							if(is_destroyed_l5(49)='0')then
								if(coll_x_l5(49)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(49)<='1';
								end if;
								if(coll_y_l5(49)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(49)<='1';
								end if;
							end if;
							if(is_destroyed_l5(48)='0')then
								if(coll_x_l5(48)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(48)<='1';
								end if;
								if(coll_y_l5(48)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(48)<='1';
								end if;
							end if;
							
							if(is_destroyed_l5(47)='0')then
								if(coll_x_l5(47)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(47)<='1';
								end if;
								if(coll_y_l5(47)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(47)<='1';
								end if;
							end if;
							if(is_destroyed_l5(46)='0')then
								if(coll_x_l5(46)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(46)<='1';
								end if;
								if(coll_y_l5(46)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(46)<='1';
								end if;
							end if;
							if(is_destroyed_l5(45)='0')then
								if(coll_x_l5(45)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(45)<='1';
								end if;
								if(coll_y_l5(45)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(45)<='1';
								end if;
							end if;						
							if(is_destroyed_l5(44)='0')then
								if(coll_x_l5(44)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(44)<='1';
								end if;
								if(coll_y_l5(44)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(44)<='1';
								end if;
							end if;						
							if(is_destroyed_l5(43)='0')then
								if(coll_x_l5(43)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(43)<='1';
								end if;
								if(coll_y_l5(43)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(43)<='1';
								end if;
							end if;
							if(is_destroyed_l5(42)='0')then
								if(coll_x_l5(42)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(42)<='1';
								end if;
								if(coll_y_l5(42)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(42)<='1';
								end if;
							end if;
							if(is_destroyed_l5(41)='0')then
								if(coll_x_l5(41)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(41)<='1';
								end if;
								if(coll_y_l5(41)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(41)<='1';
								end if;
							end if;
							if(is_destroyed_l5(40)='0')then
								if(coll_x_l5(40)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(40)<='1';
								end if;
								if(coll_y_l5(40)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(40)<='1';
								end if;
							end if;
							
							if(is_destroyed_l5(39)='0')then
								if(coll_x_l5(39)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(39)<='1';
								end if;
								if(coll_y_l5(39)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(39)<='1';
								end if;
							end if;
							if(is_destroyed_l5(38)='0')then
								if(coll_x_l5(38)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(38)<='1';
								end if;
								if(coll_y_l5(38)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(38)<='1';
								end if;
							end if;
							if(is_destroyed_l5(37)='0')then
								if(coll_x_l5(37)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(37)<='1';
								end if;
								if(coll_y_l5(37)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(37)<='1';
								end if;
							end if;						
							if(is_destroyed_l5(36)='0')then
								if(coll_x_l5(36)='1')then
									ball_x_vel<=not ball_x_vel;
									is_destroyed_l5(36)<='1';
								end if;
								if(coll_y_l5(36)='1')then
									ball_y_vel<=not ball_y_vel;
									is_destroyed_l5(36)<='1';
								end if;
							end if;


							if(ball_y>480 and isalive/=0) then--respawn ball 
								ball_x<=rand_x;
								ball_x_vel<=ball_x_vel_rand;
								bat_x<=rand_x-25;
							elsif(ball_x_vel='1' and notstarted='0' and pause='0' and stopball='0') then
								ball_x <= ball_x + 3;--move ball right
							elsif(ball_x_vel='0' and notstarted='0' and pause='0' and stopball='0') then
								ball_x <= ball_x - 3;--move ball left
							else 
								null;
							end if;

							if(ball_y>480 and isalive/=0) then--respawn ball and decrement lives
								ball_y<=450;
								ball_y_vel<='0';
								bat_y<=460;
								isalive<=isalive-1;
							elsif(ball_y_vel='1' and notstarted='0' and pause='0' and stopball='0') then
								ball_y <= ball_y + 1;--move ball down 
							elsif(ball_y_vel='0' and notstarted='0' and pause='0' and stopball='0') then
								ball_y <= ball_y - 1;--move ball up
							else
								null;
							end if;
						
							if(r_shift='0' and bat_x<590 and pause='0' and stopball='0' and ball_y<470) then
								bat_x<=bat_x+3;--move bat right
							elsif(l_shift='0' and bat_x>3 and pause='0' and stopball='0' and ball_y<470) then
								bat_x<=bat_x-3;--move bat left
							else
								null;
							end if;
							
						end if;
					end if;
							
					if(hpos>7 and hpos<104) then
						hsync<='0';	--generate the horizontal sync
					else
						hsync<='1';
					end if;
					
					if(vpos>2 and vpos<5) then
						vsync<='0';		--generate vertical sync
					else
						vsync<='1';
					end if;
			end if;
		end process;
end sync_arch;